`include "madgwickDefines.vh"

`define NUM_ELEMENTS 5000

parameter logic signed [`ACC_WIDTH-1:0] AX_TEST_VECTOR[`NUM_ELEMENTS] = {
    17'b11110111000010100,
    17'b11110110011110110,
    17'b11110101100110011,
    17'b11110100001111011,
    17'b11110011000111101,
    17'b11110010000000000,
    17'b11110001011100001,
    17'b11110000111000011,
    17'b11110000011110110,
    17'b11110000010100100,
    17'b11110000001010010,
    17'b11110000011001101,
    17'b11110000101001000,
    17'b11110000111000011,
    17'b11110000101110001,
    17'b11110000111000011,
    17'b11110001000010100,
    17'b11110001011100001,
    17'b11110001100110011,
    17'b11110001100110011,
    17'b11110001010111000,
    17'b11110000010100100,
    17'b11101111101011100,
    17'b11101110101110001,
    17'b11101101111010111,
    17'b11101100011001101,
    17'b11101011001100110,
    17'b11101001110101110,
    17'b11101000011110110,
    17'b11100110111000011,
    17'b11100101111010111,
    17'b11100110000101001,
    17'b11100110000000000,
    17'b11101001000010100,
    17'b11101100001010010,
    17'b11101011000010100,
    17'b11100100101001000,
    17'b11011110101110001,
    17'b11011001001100110,
    17'b11010101010111000,
    17'b11010101000010100,
    17'b11010111000111101,
    17'b11011001100001010,
    17'b11011011000010100,
    17'b11011100001111011,
    17'b11011100011001101,
    17'b11011100101001000,
    17'b11011100111000011,
    17'b11011101000111101,
    17'b11011101000111101,
    17'b11011101000010100,
    17'b11011101001100110,
    17'b11011101000111101,
    17'b11011101010001111,
    17'b11011101000010100,
    17'b11011101000010100,
    17'b11011100111000011,
    17'b11011100110011010,
    17'b11011100101110001,
    17'b11011100001010010,
    17'b11011011110101110,
    17'b11011011010001111,
    17'b11011011001100110,
    17'b11011010011001101,
    17'b11011000000101001,
    17'b11010101100001010,
    17'b11010100110011010,
    17'b11010110000000000,
    17'b11010111010111000,
    17'b11011001010111000,
    17'b11011011100001010,
    17'b11011110111000011,
    17'b11100001000010100,
    17'b11100010101001000,
    17'b11100010111000011,
    17'b11011101100001010,
    17'b11010100001010010,
    17'b11001110011110110,
    17'b11001011100001010,
    17'b11001010100011111,
    17'b11010000100011111,
    17'b11011101010111000,
    17'b11101101101011100,
    17'b11111010011110110,
    17'b00000001010111000,
    17'b11110100110011010,
    17'b11100100001111011,
    17'b11010111100110011,
    17'b11010000011001101,
    17'b11001110110011010,
    17'b11010010000101001,
    17'b11010110101001000,
    17'b11011010011001101,
    17'b11011100011110110,
    17'b11011100011110110,
    17'b11011010011110110,
    17'b11010111001100110,
    17'b11010000111000011,
    17'b11001011001100110,
    17'b11000110000101001,
    17'b11000100010100100,
    17'b11000101010001111,
    17'b11000011010111000,
    17'b11000100101001000,
    17'b11000111100110011,
    17'b11001011111010111,
    17'b11011000001111011,
    17'b11011111100001010,
    17'b11100100001111011,
    17'b11101000011110110,
    17'b11101001010111000,
    17'b11100011010111000,
    17'b11011101001100110,
    17'b11011000110011010,
    17'b11010111011100001,
    17'b11011000000000000,
    17'b11011000101110001,
    17'b11011000110011010,
    17'b11011000101110001,
    17'b11011000011110110,
    17'b11011000100011111,
    17'b11010111100001010,
    17'b11010111100110011,
    17'b11011000011110110,
    17'b11011000110011010,
    17'b11011010101001000,
    17'b11011011111010111,
    17'b11011100101001000,
    17'b11011101100001010,
    17'b11011110100011111,
    17'b11011111101011100,
    17'b11100000100011111,
    17'b11100010000000000,
    17'b11100010101001000,
    17'b11100011100110011,
    17'b11100011010111000,
    17'b11100000011110110,
    17'b11011011010111000,
    17'b11011001000010100,
    17'b11011010011001101,
    17'b11011011000010100,
    17'b11011010101001000,
    17'b11011010010100100,
    17'b11011010011110110,
    17'b11011000011110110,
    17'b11011010011110110,
    17'b11010101010111000,
    17'b11001100001010010,
    17'b11010110111101100,
    17'b11100000110011010,
    17'b11100000011110110,
    17'b11011111001100110,
    17'b11100101101011100,
    17'b11011100101001000,
    17'b11011101000111101,
    17'b11010110010100100,
    17'b11010010001111011,
    17'b11010011010111000,
    17'b11010110110011010,
    17'b11011001100110011,
    17'b11011011011100001,
    17'b11011100000000000,
    17'b11011010110011010,
    17'b11011001101011100,
    17'b11011001110000101,
    17'b11011100010100100,
    17'b11011111001100110,
    17'b11011101011100001,
    17'b11010111011100001,
    17'b11010100001111011,
    17'b11010010111101100,
    17'b11010011110101110,
    17'b11010101100001010,
    17'b11010110001111011,
    17'b11010110111000011,
    17'b11011000111000011,
    17'b11100001000111101,
    17'b11011110111101100,
    17'b11011011010001111,
    17'b11010110010100100,
    17'b11010111010001111,
    17'b11011001110101110,
    17'b11011001001100110,
    17'b11011111101011100,
    17'b11100110101110001,
    17'b11101000011001101,
    17'b11100001100110011,
    17'b11011001010001111,
    17'b11010100011001101,
    17'b11010100111101100,
    17'b11011000001010010,
    17'b11011100010100100,
    17'b11100001001100110,
    17'b11100010011110110,
    17'b11011111111010111,
    17'b11011011100001010,
    17'b11010101111010111,
    17'b11010011011100001,
    17'b11010010010100100,
    17'b11010001110101110,
    17'b11010011010001111,
    17'b11010111010001111,
    17'b11010110110011010,
    17'b11010101000111101,
    17'b11010111100001010,
    17'b11010111111010111,
    17'b11010110101001000,
    17'b11010111100001010,
    17'b11011011010001111,
    17'b11011101001100110,
    17'b11011101110101110,
    17'b11011100100011111,
    17'b11011001111010111,
    17'b11010110000101001,
    17'b11010011010111000,
    17'b11010001010001111,
    17'b11001111000111101,
    17'b11001100011110110,
    17'b11001010000101001,
    17'b11000111100001010,
    17'b11000101010001111,
    17'b11000100000101001,
    17'b11000101010001111,
    17'b11000111111010111,
    17'b11001011011100001,
    17'b11001110101110001,
    17'b11010010101001000,
    17'b11010100001111011,
    17'b11010101000010100,
    17'b11010100111000011,
    17'b11010100010100100,
    17'b11010100001010010,
    17'b11010100001010010,
    17'b11010100011001101,
    17'b11010100000000000,
    17'b11010010111101100,
    17'b11010001010001111,
    17'b11001110111101100,
    17'b11001101010001111,
    17'b11001100001010010,
    17'b11001011100110011,
    17'b11001011100001010,
    17'b11001011011100001,
    17'b11001011000010100,
    17'b11001010000101001,
    17'b11000100101110001,
    17'b10111111110101110,
    17'b10101010010100100,
    17'b10001111100110011,
    17'b10011001100001010,
    17'b10100110001111011,
    17'b10101110001111011,
    17'b10110100000101001,
    17'b10111101000111101,
    17'b11001000010100100,
    17'b11001100000000000,
    17'b11010000111101100,
    17'b11010100111101100,
    17'b11011010101110001,
    17'b11011110001010010,
    17'b11100000011001101,
    17'b11011111010001111,
    17'b11011100001111011,
    17'b11011001110101110,
    17'b11010110000101001,
    17'b11010010011110110,
    17'b11001110111101100,
    17'b11001100011001101,
    17'b11001001111010111,
    17'b11001000011110110,
    17'b11000110111101100,
    17'b11000111010001111,
    17'b11001000100011111,
    17'b11001010111000011,
    17'b11001101111010111,
    17'b11010010100011111,
    17'b11010101110101110,
    17'b11010111110101110,
    17'b11011010111000011,
    17'b11011110000101001,
    17'b11100000010100100,
    17'b11100010100011111,
    17'b11100010000101001,
    17'b11011101100001010,
    17'b11011010101110001,
    17'b11011001000010100,
    17'b11010111000010100,
    17'b11010100000000000,
    17'b11010001101011100,
    17'b11010000111101100,
    17'b11010000110011010,
    17'b11010000111101100,
    17'b11010001011100001,
    17'b11010000100011111,
    17'b11010000011001101,
    17'b11010000010100100,
    17'b11010000110011010,
    17'b11010001000010100,
    17'b11010001001100110,
    17'b11010001001100110,
    17'b11010001100001010,
    17'b11010001100001010,
    17'b11010001101011100,
    17'b11010010000000000,
    17'b11010010001111011,
    17'b11010010011110110,
    17'b11010010100011111,
    17'b11010010101001000,
    17'b11010010010100100,
    17'b11010010001111011,
    17'b11010010001010010,
    17'b11010010000000000,
    17'b11010001110101110,
    17'b11010001101011100,
    17'b11010001011100001,
    17'b11010001010001111,
    17'b11010001000111101,
    17'b11010001000010100,
    17'b11010001000010100,
    17'b11010000111101100,
    17'b11010001000010100,
    17'b11010001000111101,
    17'b11010001000010100,
    17'b11010001010111000,
    17'b11010001100001010,
    17'b11010001111010111,
    17'b11010010000000000,
    17'b11010010001111011,
    17'b11010010001111011,
    17'b11010010010100100,
    17'b11010010001010010,
    17'b11010010000101001,
    17'b11010010001010010,
    17'b11010010000101001,
    17'b11010010000000000,
    17'b11010001110101110,
    17'b11010001111010111,
    17'b11010001101011100,
    17'b11010001100110011,
    17'b11010001101011100,
    17'b11010001101011100,
    17'b11010001100110011,
    17'b11010001100001010,
    17'b11010001100110011,
    17'b11010001011100001,
    17'b11010001101011100,
    17'b11010001101011100,
    17'b11010001110000101,
    17'b11010001110101110,
    17'b11010001111010111,
    17'b11010010000000000,
    17'b11010010001010010,
    17'b11010010001111011,
    17'b11010010001010010,
    17'b11010010001111011,
    17'b11010010001111011,
    17'b11010010010100100,
    17'b11010010000101001,
    17'b11010010001010010,
    17'b11010010000101001,
    17'b11010001111010111,
    17'b11010001111010111,
    17'b11010001110101110,
    17'b11010001111010111,
    17'b11010001111010111,
    17'b11010100111101100,
    17'b11010111110000101,
    17'b11011000001010010,
    17'b11010100100011111,
    17'b11010011100001010,
    17'b11010011010111000,
    17'b11010011000010100,
    17'b11010011001100110,
    17'b11010010000101001,
    17'b11010000011110110,
    17'b11001110101110001,
    17'b11001011100001010,
    17'b11001011101011100,
    17'b11001100001010010,
    17'b11001101001100110,
    17'b11010001000010100,
    17'b11010010001010010,
    17'b11010010010100100,
    17'b11010001111010111,
    17'b11010000101110001,
    17'b11010000011110110,
    17'b11010000100011111,
    17'b11010001010001111,
    17'b11010010010100100,
    17'b11010011000111101,
    17'b11010011011100001,
    17'b11010011001100110,
    17'b11010010110011010,
    17'b11010010001010010,
    17'b11010010100011111,
    17'b11010010111000011,
    17'b11010011000111101,
    17'b11010010111000011,
    17'b11010010011001101,
    17'b11010010000000000,
    17'b11010001010111000,
    17'b11010001010111000,
    17'b11010001010111000,
    17'b11010001101011100,
    17'b11010010000000000,
    17'b10111100101110001,
    17'b10111010000101001,
    17'b11001000100011111,
    17'b11011011101011100,
    17'b11001011001100110,
    17'b11001011100001010,
    17'b10111101100001010,
    17'b10110111110101110,
    17'b10111011100001010,
    17'b11000000000101001,
    17'b11000100111000011,
    17'b11001000010100100,
    17'b11001100010100100,
    17'b11001110110011010,
    17'b11001110101001000,
    17'b11001110010100100,
    17'b11001110110011010,
    17'b11010001011100001,
    17'b11010110000000000,
    17'b11000111101011100,
    17'b11100101101011100,
    17'b00001001010001111,
    17'b00010001110000101,
    17'b00010010000101001,
    17'b00010001100110011,
    17'b00010000011110110,
    17'b00001011000010100,
    17'b11111011000111101,
    17'b11100111000111101,
    17'b11010101000111101,
    17'b10111110011001101,
    17'b10101000010100100,
    17'b10011010001111011,
    17'b10001111110000101,
    17'b10000111110101110,
    17'b10000101000010100,
    17'b10001000011001101,
    17'b10001100011110110,
    17'b10010100000101001,
    17'b10100000100011111,
    17'b10101100011110110,
    17'b10111001001100110,
    17'b11001011010111000,
    17'b11010101011100001,
    17'b11011110000101001,
    17'b11100100011001101,
    17'b11101010111000011,
    17'b11101111010001111,
    17'b11110011000010100,
    17'b11110110011110110,
    17'b11111000101001000,
    17'b11110111011100001,
    17'b11110000001010010,
    17'b11101100001010010,
    17'b11100111010001111,
    17'b11100000000101001,
    17'b11011110000000000,
    17'b11011100010100100,
    17'b11011001011100001,
    17'b11010100010100100,
    17'b11010000010100100,
    17'b11001100011110110,
    17'b11001011100001010,
    17'b11001101000010100,
    17'b11001110000000000,
    17'b11001110101001000,
    17'b11001111000010100,
    17'b11001110001111011,
    17'b11001101010001111,
    17'b11001100011110110,
    17'b11001011100110011,
    17'b11010000111101100,
    17'b11010011010001111,
    17'b11010011101011100,
    17'b11010100000000000,
    17'b11010011000010100,
    17'b11010000011110110,
    17'b11001111110000101,
    17'b11010000000000000,
    17'b11010001000111101,
    17'b11010010011110110,
    17'b11010010011001101,
    17'b11010010000101001,
    17'b11010001111010111,
    17'b11010001000010100,
    17'b11010000111101100,
    17'b11010001000010100,
    17'b11010010000000000,
    17'b11010010101110001,
    17'b11010011100001010,
    17'b11010100000101001,
    17'b11010100011001101,
    17'b11010100111000011,
    17'b11010100111000011,
    17'b11010101001100110,
    17'b11010101001100110,
    17'b11010101010111000,
    17'b11010101000111101,
    17'b11010100010100100,
    17'b11010011101011100,
    17'b11010010101110001,
    17'b11010010001010010,
    17'b11010011010001111,
    17'b11010011110000101,
    17'b11010001010001111,
    17'b11001111111010111,
    17'b11010000000101001,
    17'b11001101000111101,
    17'b11001100111000011,
    17'b11001101100001010,
    17'b11100111111010111,
    17'b00100000110011010,
    17'b00000010011001101,
    17'b11010010010100100,
    17'b11001011100110011,
    17'b11000011001100110,
    17'b11010001000010100,
    17'b11001001111010111,
    17'b11000000011110110,
    17'b10111100110011010,
    17'b11000111000111101,
    17'b11010000011001101,
    17'b11010001000111101,
    17'b11010101010001111,
    17'b11010100100011111,
    17'b11001101010001111,
    17'b11000110001111011,
    17'b11000011111010111,
    17'b11000001101011100,
    17'b11000100110011010,
    17'b11001000100011111,
    17'b11001001110101110,
    17'b11001111110000101,
    17'b11011101100001010,
    17'b11101100111101100,
    17'b11101110100011111,
    17'b11011000011110110,
    17'b11000010000000000,
    17'b10110000100011111,
    17'b10101001110000101,
    17'b10110001100001010,
    17'b10111100000000000,
    17'b11000100100011111,
    17'b11001000001010010,
    17'b11000110111101100,
    17'b11000011101011100,
    17'b11000010000000000,
    17'b11000010011110110,
    17'b11000011110000101,
    17'b11000011101011100,
    17'b11000010000101001,
    17'b11000010001111011,
    17'b11000100000101001,
    17'b11000101110101110,
    17'b11000111110000101,
    17'b11001001000010100,
    17'b11001001101011100,
    17'b11001001101011100,
    17'b11001000111101100,
    17'b11001001010111000,
    17'b11001010100011111,
    17'b11001010111101100,
    17'b11001010100011111,
    17'b11001010001010010,
    17'b11001001101011100,
    17'b11000111110101110,
    17'b11000100011001101,
    17'b11000000001010010,
    17'b10111101000010100,
    17'b10111011001100110,
    17'b10111010001111011,
    17'b10111001001100110,
    17'b10111000000000000,
    17'b10110111101011100,
    17'b10111000001010010,
    17'b10111001000010100,
    17'b10111011000010100,
    17'b10111101000111101,
    17'b10111111000111101,
    17'b11000000111101100,
    17'b11000010100011111,
    17'b11000110101110001,
    17'b11001001000111101,
    17'b11001010101110001,
    17'b11001100011001101,
    17'b11001110100011111,
    17'b11001000011110110,
    17'b11000100011110110,
    17'b11000111110101110,
    17'b11010000000101001,
    17'b11010111010001111,
    17'b11011100011110110,
    17'b11011111010001111,
    17'b11100000011110110,
    17'b11100000111000011,
    17'b11100011010111000,
    17'b11100100111101100,
    17'b11100110001010010,
    17'b11101001010111000,
    17'b11101010111000011,
    17'b11101000111101100,
    17'b11101010101110001,
    17'b11101010101110001,
    17'b11101011010111000,
    17'b11101100100011111,
    17'b11101011110101110,
    17'b11101010110011010,
    17'b11101010001111011,
    17'b11101000100011111,
    17'b11101001010001111,
    17'b11101001000010100,
    17'b11101001110101110,
    17'b11101000000101001,
    17'b11101000001010010,
    17'b11100111110101110,
    17'b11100100000000000,
    17'b11100011010001111,
    17'b11100101101011100,
    17'b11100111010111000,
    17'b11101010001111011,
    17'b11100101010111000,
    17'b11100001011100001,
    17'b11011110011110110,
    17'b11100011010001111,
    17'b00001000011110110,
    17'b00111100100011111,
    17'b01001111010001111,
    17'b00110111000010100,
    17'b00100100111000011,
    17'b00011010110011010,
    17'b00010011000010100,
    17'b00000011110101110,
    17'b00000000001010010,
    17'b00001001100110011,
    17'b00010111010111000,
    17'b00100000001111011,
    17'b00100101000010100,
    17'b00100111111010111,
    17'b00101000000000000,
    17'b00100011111010111,
    17'b00011101100001010,
    17'b00011011011100001,
    17'b00011010000000000,
    17'b00010111001100110,
    17'b00010011000111101,
    17'b00010001100110011,
    17'b00010010000101001,
    17'b00010010010100100,
    17'b00010010000101001,
    17'b00010011000111101,
    17'b00001111111010111,
    17'b00001001101011100,
    17'b11111110100011111,
    17'b11110001111010111,
    17'b11101110111000011,
    17'b11110100011001101,
    17'b11111010001010010,
    17'b00000001110101110,
    17'b00001011100001010,
    17'b00001110000000000,
    17'b00001110011110110,
    17'b00010000000101001,
    17'b00010010011001101,
    17'b00010100001010010,
    17'b00010100001111011,
    17'b00010001010001111,
    17'b00001110001111011,
    17'b00001110000101001,
    17'b00010000011110110,
    17'b00010010110011010,
    17'b00010100011110110,
    17'b00010101111010111,
    17'b00010110011001101,
    17'b00010110001010010,
    17'b00010100011001101,
    17'b00010100110011010,
    17'b00011000111000011,
    17'b00100010000101001,
    17'b00101011111010111,
    17'b00110001001100110,
    17'b00110111000111101,
    17'b00111000111101100,
    17'b00111011101011100,
    17'b00111100101001000,
    17'b00111000011110110,
    17'b00110011011100001,
    17'b00101110011001101,
    17'b00101000101110001,
    17'b00100000001010010,
    17'b00011101110101110,
    17'b00011111010111000,
    17'b00100010111000011,
    17'b00100110100011111,
    17'b00101000000101001,
    17'b00101000110011010,
    17'b00101001101011100,
    17'b00101010100011111,
    17'b00101010101110001,
    17'b00101001110101110,
    17'b00101000000101001,
    17'b00100110001111011,
    17'b00100011010001111,
    17'b00100001000111101,
    17'b00011110111101100,
    17'b00011101000010100,
    17'b00011100101110001,
    17'b00011101100001010,
    17'b00011110011110110,
    17'b00011110110011010,
    17'b00011110101110001,
    17'b00011110010100100,
    17'b00011111111010111,
    17'b00011101111010111,
    17'b00011111010001111,
    17'b00011110111101100,
    17'b00100001010001111,
    17'b00100011000111101,
    17'b00100011100110011,
    17'b00100001011100001,
    17'b00100010011110110,
    17'b00100001000010100,
    17'b00100000101001000,
    17'b00100001100110011,
    17'b00100000000101001,
    17'b00011100010100100,
    17'b00011000111000011,
    17'b00010100111000011,
    17'b00100111000111101,
    17'b00010101000111101,
    17'b00000100000000000,
    17'b00000110000101001,
    17'b00001011000111101,
    17'b00000001010111000,
    17'b11111010110011010,
    17'b00000111000111101,
    17'b00010110000101001,
    17'b00010010101001000,
    17'b00001101000010100,
    17'b00000111110000101,
    17'b00000011001100110,
    17'b11111111101011100,
    17'b11111111110101110,
    17'b00000001000111101,
    17'b00000010011110110,
    17'b00000010100011111,
    17'b00000010111101100,
    17'b00000011100110011,
    17'b00000100100011111,
    17'b00000101010111000,
    17'b00000110000101001,
    17'b00000110100011111,
    17'b00000110111101100,
    17'b00001001111010111,
    17'b00001011100110011,
    17'b00001100111101100,
    17'b00001111110101110,
    17'b00010011000010100,
    17'b00010100000000000,
    17'b00010101010001111,
    17'b00011001000010100,
    17'b00011001011100001,
    17'b00011011111010111,
    17'b00011100001111011,
    17'b00011110100011111,
    17'b00011110110011010,
    17'b00011111100001010,
    17'b00100000000000000,
    17'b00011111110101110,
    17'b00011111110000101,
    17'b00011111000111101,
    17'b00011111111010111,
    17'b00011111110000101,
    17'b00011110011001101,
    17'b00011010111101100,
    17'b00010101111010111,
    17'b00010010001010010,
    17'b00001101101011100,
    17'b00001001100110011,
    17'b00000111110000101,
    17'b00000101000111101,
    17'b00000101111010111,
    17'b00000100110011010,
    17'b00000010101001000,
    17'b00000110101001000,
    17'b00001011101011100,
    17'b00001101001100110,
    17'b00001101000010100,
    17'b00001110001010010,
    17'b00010000000101001,
    17'b00010010000101001,
    17'b00010011000010100,
    17'b00010100010100100,
    17'b00010110000101001,
    17'b00010111110101110,
    17'b00011001100001010,
    17'b00011010011001101,
    17'b00011100001111011,
    17'b00011101101011100,
    17'b00011111001100110,
    17'b00100000111101100,
    17'b00100011000111101,
    17'b00100100101001000,
    17'b00100101110000101,
    17'b00100101111010111,
    17'b00100110011001101,
    17'b00100110000000000,
    17'b00100100100011111,
    17'b00100010110011010,
    17'b00100001011100001,
    17'b00011100101110001,
    17'b00011101110000101,
    17'b00011011111010111,
    17'b00011000100011111,
    17'b00010110010100100,
    17'b00011001110000101,
    17'b00010100000000000,
    17'b00010110000000000,
    17'b00011000000000000,
    17'b00010111010111000,
    17'b00010110011001101,
    17'b00010101001100110,
    17'b00010100011001101,
    17'b00010010100011111,
    17'b00010001101011100,
    17'b00010001111010111,
    17'b00010001100001010,
    17'b00010001100001010,
    17'b00010000101110001,
    17'b00001111110101110,
    17'b00001110101001000,
    17'b00001111000010100,
    17'b00001101110101110,
    17'b00001101000111101,
    17'b00001100011001101,
    17'b00001100000101001,
    17'b00001011010001111,
    17'b00001010101001000,
    17'b00001001000010100,
    17'b00000111101011100,
    17'b00000110101001000,
    17'b00000100010100100,
    17'b00000011100110011,
    17'b00000010111101100,
    17'b00000010001111011,
    17'b00000001100110011,
    17'b00000001100001010,
    17'b00000001011100001,
    17'b00000001010111000,
    17'b00000001110000101,
    17'b00000010000101001,
    17'b00000010011001101,
    17'b00000010101110001,
    17'b00000011100110011,
    17'b00000011111010111,
    17'b00000100000000000,
    17'b00000011110000101,
    17'b00000010111000011,
    17'b00000010011001101,
    17'b00000001110000101,
    17'b00000001000010100,
    17'b00000000001010010,
    17'b11111111000010100,
    17'b11111110001010010,
    17'b11111101010111000,
    17'b11111101000010100,
    17'b11111100100011111,
    17'b11111100011001101,
    17'b11111100000000000,
    17'b11111100001010010,
    17'b11111100000000000,
    17'b11111100111000011,
    17'b11111110010100100,
    17'b11111111100001010,
    17'b00000000000101001,
    17'b00000000011001101,
    17'b00000001000010100,
    17'b00000010000101001,
    17'b00000001100001010,
    17'b11111111111010111,
    17'b11111110110011010,
    17'b11111110101110001,
    17'b11111110010100100,
    17'b11111101010001111,
    17'b11111100101001000,
    17'b11111011000111101,
    17'b11111011100001010,
    17'b11111010101110001,
    17'b11111010010100100,
    17'b11111000110011010,
    17'b11110111010001111,
    17'b11110010100011111,
    17'b11110100101110001,
    17'b11110101010111000,
    17'b11110100100011111,
    17'b11110101100001010,
    17'b11110110010100100,
    17'b11110111011100001,
    17'b11110110001111011,
    17'b11110111000111101,
    17'b11111011000010100,
    17'b11111011010111000,
    17'b11111010110011010,
    17'b11111000000101001,
    17'b11101001000111101,
    17'b11011001101011100,
    17'b11010001000111101,
    17'b11001111000010100,
    17'b10111100101001000,
    17'b10110001100110011,
    17'b10111100110011010,
    17'b11010011011100001,
    17'b11100110101110001,
    17'b11110101111010111,
    17'b00110001011100001,
    17'b01010100011110110,
    17'b01101000001111011,
    17'b01011010000101001,
    17'b00111001000010100,
    17'b00100010110011010,
    17'b00010011100110011,
    17'b00000101111010111,
    17'b11110011100110011,
    17'b11101101101011100,
    17'b11101111011100001,
    17'b11110101000111101,
    17'b11110001100110011,
    17'b11101011111010111,
    17'b11101000000000000,
    17'b11101110011110110,
    17'b11111110111000011,
    17'b00000011000010100,
    17'b00000100000101001,
    17'b00000100010100100,
    17'b00000100000000000,
    17'b00010001100110011,
    17'b00010010101110001,
    17'b00001001010001111,
    17'b11111101110101110,
    17'b11111001110101110,
    17'b11110111000111101,
    17'b11111000011110110,
    17'b11111011100110011,
    17'b11111111101011100,
    17'b11110111000010100,
    17'b11101100111000011,
    17'b11110000001111011,
    17'b11101111010001111,
    17'b11101100110011010,
    17'b11101011010111000,
    17'b11101101110000101,
    17'b11110101000111101,
    17'b11110101100001010,
    17'b11101100100011111,
    17'b11101111011100001,
    17'b11110100101001000,
    17'b11110110110011010,
    17'b11111000111101100,
    17'b11111110001010010,
    17'b00001000101110001,
    17'b00011000101110001,
    17'b00101110101001000,
    17'b00110100000101001,
    17'b00101010011110110,
    17'b00100000101110001,
    17'b00011110111101100,
    17'b00100111101011100,
    17'b00100100000101001,
    17'b00100011001100110,
    17'b00011010111101100,
    17'b00101011000010100,
    17'b00100101011100001,
    17'b01010000100011111,
    17'b00111110100011111,
    17'b00110010101110001,
    17'b00101111111010111,
    17'b00101100011001101,
    17'b00110000000101001,
    17'b00110011110101110,
    17'b00110001010111000,
    17'b00110000111101100,
    17'b00101100011001101,
    17'b00101000110011010,
    17'b00100110110011010,
    17'b00100110110011010,
    17'b00100110010100100,
    17'b00100110111101100,
    17'b00100111000111101,
    17'b00100110010100100,
    17'b00101000101001000,
    17'b00101010100011111,
    17'b00110100000101001,
    17'b00111010010100100,
    17'b01000001110000101,
    17'b01001001011100001,
    17'b01010000110011010,
    17'b01011000111101100,
    17'b01011101010001111,
    17'b01011110110011010,
    17'b01011100110011010,
    17'b01010101100110011,
    17'b01001110101001000,
    17'b01000111110101110,
    17'b01000001101011100,
    17'b00111011110000101,
    17'b00110111111010111,
    17'b00110100101001000,
    17'b00110001110101110,
    17'b00101110110011010,
    17'b00101101011100001,
    17'b00101101010111000,
    17'b00110000000000000,
    17'b00110100101110001,
    17'b00110111010111000,
    17'b00111011000010100,
    17'b00111110011110110,
    17'b01000000111000011,
    17'b01000010111101100,
    17'b01000100110011010,
    17'b01000111100001010,
    17'b01001011010111000,
    17'b01001111010111000,
    17'b01010000110011010,
    17'b01010001101011100,
    17'b01010001001100110,
    17'b01001111010001111,
    17'b01001100011001101,
    17'b01000111100110011,
    17'b01000011110000101,
    17'b01000000100011111,
    17'b00111110000000000,
    17'b00111001010001111,
    17'b00110111110000101,
    17'b00110111110101110,
    17'b00110110110011010,
    17'b00111011000111101,
    17'b00111110111000011,
    17'b01000001010111000,
    17'b01000011111010111,
    17'b01001110011001101,
    17'b01010011011100001,
    17'b01010111100110011,
    17'b01011001110000101,
    17'b01011101110101110,
    17'b01011000100011111,
    17'b01011111111010111,
    17'b01011110111101100,
    17'b01011100000101001,
    17'b01011011000010100,
    17'b01010101110000101,
    17'b01001111010111000,
    17'b01001000011110110,
    17'b01000111100110011,
    17'b01000111000111101,
    17'b01000111111010111,
    17'b01001011011100001,
    17'b01001111110101110,
    17'b01010011100110011,
    17'b01010110011110110,
    17'b01010110100011111,
    17'b01010100101110001,
    17'b01010001101011100,
    17'b01001100000000000,
    17'b01000110000101001,
    17'b00111110011110110,
    17'b00110110101110001,
    17'b00101110011001101,
    17'b00101010000101001,
    17'b00100111000111101,
    17'b00100111110101110,
    17'b00100100101001000,
    17'b00011101111010111,
    17'b00011010101001000,
    17'b00011001010111000,
    17'b00011001110101110,
    17'b00011011011100001,
    17'b00011110001010010,
    17'b00100001000111101,
    17'b00100010110011010,
    17'b00100010001010010,
    17'b00011111100001010,
    17'b00011100111101100,
    17'b00011010100011111,
    17'b00011001010111000,
    17'b00011001010111000,
    17'b00011011000010100,
    17'b00011100101110001,
    17'b00011100100011111,
    17'b00010010101001000,
    17'b00000101111010111,
    17'b00001100101110001,
    17'b00001001001100110,
    17'b11111100000101001,
    17'b11110001110101110,
    17'b11101110010100100,
    17'b11101100000101001,
    17'b11100111101011100,
    17'b11100010101001000,
    17'b11011110001111011,
    17'b11011100010100100,
    17'b11011100001010010,
    17'b11011000011001101,
    17'b11010001110000101,
    17'b11010100101001000,
    17'b11010100000000000,
    17'b11010011001100110,
    17'b11011001110000101,
    17'b11011110101001000,
    17'b11011001100110011,
    17'b11010111010111000,
    17'b11011001001100110,
    17'b11011101100001010,
    17'b11100001000111101,
    17'b11100000000101001,
    17'b11011110101001000,
    17'b11011100111101100,
    17'b11010100110011010,
    17'b11001110001010010,
    17'b11010100111101100,
    17'b11010111110000101,
    17'b11011011001100110,
    17'b11100000100011111,
    17'b11100000001111011,
    17'b11011011001100110,
    17'b11010111011100001,
    17'b11010100111101100,
    17'b11010011101011100,
    17'b11010001110101110,
    17'b11010000001111011,
    17'b11001110001111011,
    17'b11001100011001101,
    17'b11001010011110110,
    17'b11001011001100110,
    17'b11001100101110001,
    17'b11001110001010010,
    17'b11001111010111000,
    17'b11001111101011100,
    17'b11010011110000101,
    17'b11010110100011111,
    17'b11011011000111101,
    17'b11011100111000011,
    17'b11001111110000101,
    17'b11001011110000101,
    17'b11001100111000011,
    17'b11010000111000011,
    17'b11010110000101001,
    17'b11011011101011100,
    17'b11100000011110110,
    17'b11100011011100001,
    17'b11111101110000101,
    17'b11101110110011010,
    17'b11011110001111011,
    17'b11001110011001101,
    17'b11001011010001111,
    17'b11000110011110110,
    17'b11000111100110011,
    17'b11001111000010100,
    17'b11010100100011111,
    17'b11011000100011111,
    17'b11011010111101100,
    17'b11011011111010111,
    17'b11011010001010010,
    17'b11010110001010010,
    17'b11010001101011100,
    17'b11000100110011010,
    17'b11000110100011111,
    17'b11001011000010100,
    17'b11010010011110110,
    17'b11010111011100001,
    17'b11010101011100001,
    17'b11001111010001111,
    17'b11010000000101001,
    17'b11010001101011100,
    17'b11010001010111000,
    17'b11010001000111101,
    17'b11010000101110001,
    17'b11010010011110110,
    17'b11010011010111000,
    17'b11010000010100100,
    17'b11001110111000011,
    17'b11001110011110110,
    17'b11001101001100110,
    17'b11001100000000000,
    17'b11001101100001010,
    17'b11010010010100100,
    17'b11011001101011100,
    17'b11011101110101110,
    17'b11100000110011010,
    17'b11100010110011010,
    17'b11100100001010010,
    17'b11100011101011100,
    17'b11011110000000000,
    17'b11001010000000000,
    17'b10111001110101110,
    17'b11001000110011010,
    17'b11011011100110011,
    17'b11101010000000000,
    17'b11110100110011010,
    17'b11111101010001111,
    17'b11111110001111011,
    17'b11111111100001010,
    17'b00101100010100100,
    17'b00110100111101100,
    17'b00011001100110011,
    17'b11111101011100001,
    17'b11110011110000101,
    17'b11110101011100001,
    17'b11110110110011010,
    17'b11111001010001111,
    17'b11111111101011100,
    17'b00000100110011010,
    17'b00001001001100110,
    17'b00001100110011010,
    17'b00001111110000101,
    17'b00010010010100100,
    17'b00010110101001000,
    17'b00011111010001111,
    17'b00101001101011100,
    17'b00100110110011010,
    17'b00011111010001111,
    17'b00010110001111011,
    17'b00001111100001010,
    17'b00001111000111101,
    17'b00010010001111011,
    17'b00010110001111011,
    17'b00011011110101110,
    17'b00011110011110110,
    17'b00100000101001000,
    17'b00100010000101001,
    17'b00100011000111101,
    17'b00100100111101100,
    17'b00100110101001000,
    17'b00101000100011111,
    17'b00101010001010010,
    17'b00101100101110001,
    17'b00101110010100100,
    17'b00101111101011100,
    17'b00110001000111101,
    17'b00110100010100100,
    17'b00111000001010010,
    17'b00111100011110110,
    17'b01000000101110001,
    17'b01000011101011100,
    17'b01000101001100110,
    17'b01000101001100110,
    17'b01000101000010100,
    17'b01000101000111101,
    17'b01000101011100001,
    17'b01000101010001111,
    17'b01000100001010010,
    17'b01000011010001111,
    17'b01000001011100001,
    17'b00111111111010111,
    17'b00111110000000000,
    17'b00111100001010010,
    17'b00111011000010100,
    17'b00111010011110110,
    17'b00111011100001010,
    17'b00111101010001111,
    17'b00111111100110011,
    17'b01000010101110001,
    17'b01000110111101100,
    17'b01001010101110001,
    17'b01001010101001000,
    17'b01001010001010010,
    17'b01000111110101110,
    17'b01000101010111000,
    17'b00111110011110110,
    17'b00111110011001101,
    17'b00111111010001111,
    17'b01000000010100100,
    17'b01000001010111000,
    17'b01000001110000101,
    17'b01000010110011010,
    17'b01000011111010111,
    17'b01000101000111101,
    17'b01000110101001000,
    17'b01000111110000101,
    17'b01001000011001101,
    17'b01001001000010100,
    17'b01001001110101110,
    17'b01001011010111000,
    17'b01001101010001111,
    17'b01001110001010010,
    17'b01001101000010100,
    17'b01001011101011100,
    17'b01001001110101110,
    17'b01000111000010100,
    17'b01000100011110110,
    17'b00111110011110110,
    17'b00111001000010100,
    17'b00110111100001010,
    17'b00111010101001000,
    17'b00111111001100110,
    17'b01000010011110110,
    17'b01000011100001010,
    17'b01000010010100100,
    17'b01000000001111011,
    17'b00111110011110110,
    17'b00111101100001010,
    17'b00111110000101001,
    17'b00111111110101110,
    17'b01000010001111011,
    17'b01000110110011010,
    17'b01001001001100110,
    17'b01001010010100100,
    17'b01001011010001111,
    17'b01001100111000011,
    17'b01001101110000101,
    17'b01001110011001101,
    17'b01001110101001000,
    17'b01001110101110001,
    17'b01001110011110110,
    17'b01001110001010010,
    17'b01001110000101001,
    17'b01001101110101110,
    17'b01001101100001010,
    17'b01001100111000011,
    17'b01001011110101110,
    17'b01001010101001000,
    17'b01001001011100001,
    17'b01001001010111000,
    17'b01001001010001111,
    17'b01001000101001000,
    17'b01000111100001010,
    17'b01000110000101001,
    17'b01000101100001010,
    17'b01000100110011010,
    17'b01000100011001101,
    17'b01000100100011111,
    17'b01000101000111101,
    17'b01000100111000011,
    17'b01000101000010100,
    17'b01000100110011010,
    17'b01000100110011010,
    17'b01000101010001111,
    17'b01000101100001010,
    17'b01000110001010010,
    17'b01000111000010100,
    17'b01000111100001010,
    17'b01000111000111101,
    17'b01000110001010010,
    17'b01000011111010111,
    17'b01000000000000000,
    17'b00111111001100110,
    17'b00111111001100110,
    17'b00111001110000101,
    17'b00111000000000000,
    17'b00111101011100001,
    17'b01000100001111011,
    17'b01001011010001111,
    17'b01010001010001111,
    17'b01010011101011100,
    17'b01010101001100110,
    17'b01010101000010100,
    17'b01010110011110110,
    17'b01010110101110001,
    17'b01010001011100001,
    17'b01001100011110110,
    17'b01001000000000000,
    17'b01000011010001111,
    17'b00111110001111011,
    17'b00111011010111000,
    17'b00111001000010100,
    17'b00110111100001010,
    17'b00110110011110110,
    17'b00110110111101100,
    17'b00111000000000000,
    17'b00111001111010111,
    17'b00111101000010100,
    17'b01010110101001000,
    17'b01000101101011100,
    17'b00101101100110011,
    17'b00101000100011111,
    17'b00101110111101100,
    17'b00111110011110110,
    17'b01000111100110011,
    17'b01000001110101110,
    17'b00110110010100100,
    17'b00110011000111101,
    17'b00111010000101001,
    17'b01000011110000101,
    17'b01001011010111000,
    17'b01001011101011100,
    17'b00111101000010100,
    17'b00110100001010010,
    17'b00110011001100110,
    17'b00110111100001010,
    17'b00111010001111011,
    17'b00111100011110110,
    17'b00111101000111101,
    17'b00111100111101100,
    17'b00111100001010010,
    17'b00111011100110011,
    17'b00111010000000000,
    17'b00111000011110110,
    17'b00110111000111101,
    17'b00110100111000011,
    17'b00110001110101110,
    17'b00110000000101001,
    17'b00101110101110001,
    17'b00101011101011100,
    17'b00101000101110001,
    17'b00110101110000101,
    17'b01000110101110001,
    17'b00111001000010100,
    17'b00110000011110110,
    17'b00001111010001111,
    17'b00001101111010111,
    17'b00010100101110001,
    17'b00100000100011111,
    17'b00100110100011111,
    17'b00110111011100001,
    17'b00111101110101110,
    17'b00111011100110011,
    17'b00111000111101100,
    17'b00110011101011100,
    17'b00101011100110011,
    17'b00100111000010100,
    17'b00100000101001000,
    17'b00100000011001101,
    17'b00100001001100110,
    17'b00100001100110011,
    17'b00100010001111011,
    17'b00100011001100110,
    17'b00100011111010111,
    17'b00100010111101100,
    17'b00011110110011010,
    17'b00011011010001111,
    17'b00010111101011100,
    17'b00010101000010100,
    17'b00010001101011100,
    17'b00001111011100001,
    17'b00001110011110110,
    17'b00001110000000000,
    17'b00001101011100001,
    17'b00001101001100110,
    17'b00001100111000011,
    17'b00001101000111101,
    17'b00001101101011100,
    17'b00001110101110001,
    17'b00010000001111011,
    17'b00010010001010010,
    17'b00010011110000101,
    17'b00010100111101100,
    17'b00010101010001111,
    17'b00010110000000000,
    17'b00010110000000000,
    17'b00010100111000011,
    17'b00010011001100110,
    17'b00010010010100100,
    17'b00010001000111101,
    17'b00010000000101001,
    17'b00001110110011010,
    17'b00001101010001111,
    17'b00001011011100001,
    17'b00001000111000011,
    17'b00000111111010111,
    17'b00000111000111101,
    17'b00000110011110110,
    17'b00000101011100001,
    17'b00000100110011010,
    17'b00000011110000101,
    17'b00000011000111101,
    17'b00000010110011010,
    17'b00000011110000101,
    17'b00001001100001010,
    17'b00001000101001000,
    17'b00000111100001010,
    17'b00001000101001000,
    17'b00001001000111101,
    17'b00001001100001010,
    17'b00001100000101001,
    17'b00001110001010010,
    17'b00001001010111000,
    17'b00001000011001101,
    17'b00000111011100001,
    17'b00000110010100100,
    17'b00000101010111000,
    17'b00000011100001010,
    17'b00000100001111011,
    17'b00000101100001010,
    17'b00000101100001010,
    17'b00000011111010111,
    17'b00000011111010111,
    17'b00000000100011111,
    17'b00000010011001101,
    17'b11111111100001010,
    17'b11111100100011111,
    17'b11111010001010010,
    17'b11111000111000011,
    17'b11110101100001010,
    17'b11110011001100110,
    17'b11110010111101100,
    17'b11110101011100001,
    17'b11111001000111101,
    17'b11111110011110110,
    17'b00000010101001000,
    17'b00000101001100110,
    17'b00001100101001000,
    17'b00001010100011111,
    17'b00000101001100110,
    17'b00000000101110001,
    17'b11111100101001000,
    17'b11111001011100001,
    17'b11111001000111101,
    17'b11111001101011100,
    17'b11111010110011010,
    17'b11111100001010010,
    17'b11111101101011100,
    17'b11111101101011100,
    17'b11111100001111011,
    17'b11111000111101100,
    17'b11110100111101100,
    17'b11110000111000011,
    17'b11101111100001010,
    17'b11101111100001010,
    17'b11110000000101001,
    17'b11110001010001111,
    17'b11110011000010100,
    17'b11110100101001000,
    17'b11110110001010010,
    17'b11110111100110011,
    17'b11111001101011100,
    17'b11111100000000000,
    17'b11111010001010010,
    17'b11111000001010010,
    17'b11110111001100110,
    17'b11110011111010111,
    17'b11110011100001010,
    17'b11110011101011100,
    17'b11110010111101100,
    17'b11110010101001000,
    17'b11110011100110011,
    17'b11110101010001111,
    17'b11110101010111000,
    17'b11110100000101001,
    17'b11110011100001010,
    17'b11110011100110011,
    17'b11110110000101001,
    17'b11111001100110011,
    17'b11111011001100110,
    17'b11111001010001111,
    17'b11110111100001010,
    17'b11110101101011100,
    17'b11110100010100100,
    17'b11110011000010100,
    17'b11110011000111101,
    17'b11110010010100100,
    17'b11110001100110011,
    17'b11110001100110011,
    17'b11110001000010100,
    17'b11110000011110110,
    17'b11110000101001000,
    17'b11110010000101001,
    17'b11110011000111101,
    17'b11110100000101001,
    17'b11111000010100100,
    17'b00000110110011010,
    17'b00000101000111101,
    17'b11111101001100110,
    17'b11111001110000101,
    17'b11110111000010100,
    17'b11110011010111000,
    17'b11110001100110011,
    17'b11110001101011100,
    17'b11110010000000000,
    17'b11110010111000011,
    17'b11110100111000011,
    17'b11110111101011100,
    17'b11111001011100001,
    17'b11111010001010010,
    17'b11111010100011111,
    17'b11111011010111000,
    17'b11111011111010111,
    17'b11111100101001000,
    17'b11111101011100001,
    17'b11111101100001010,
    17'b11111100101001000,
    17'b11111100011110110,
    17'b11111011101011100,
    17'b11111010101110001,
    17'b11111001110101110,
    17'b11111001011100001,
    17'b11111001011100001,
    17'b11111001100110011,
    17'b11111011100110011,
    17'b11111101100001010,
    17'b11111111111010111,
    17'b00000010010100100,
    17'b00000101111010111,
    17'b00001000100011111,
    17'b00001010101001000,
    17'b00001100011110110,
    17'b00001110111000011,
    17'b00010000011001101,
    17'b00010001100110011,
    17'b00010011000010100,
    17'b00010100101110001,
    17'b00010110101001000,
    17'b00010111100110011,
    17'b00011000100011111,
    17'b00011001101011100,
    17'b00011010100011111,
    17'b00011010101110001,
    17'b00011010000101001,
    17'b00011001010111000,
    17'b00011000101001000,
    17'b00011000001111011,
    17'b00011000100011111,
    17'b00011010001010010,
    17'b00011100111101100,
    17'b00100001010111000,
    17'b00100101000010100,
    17'b00101000011110110,
    17'b00101011100001010,
    17'b00101101000111101,
    17'b00101101001100110,
    17'b00101011101011100,
    17'b00101001010111000,
    17'b00100111010111000,
    17'b00100101011100001,
    17'b00100011110101110,
    17'b00100001101011100,
    17'b00011111000010100,
    17'b00011110001010010,
    17'b00011110100011111,
    17'b00011100011001101,
    17'b00011001110000101,
    17'b00011000101001000,
    17'b00011001010001111,
    17'b00011011101011100,
    17'b00011110011110110,
    17'b00011111001100110,
    17'b00011110011001101,
    17'b00011100110011010,
    17'b00011011011100001,
    17'b00011010110011010,
    17'b00011010111000011,
    17'b00011010111000011,
    17'b00011011000111101,
    17'b00011011010001111,
    17'b00011011000111101,
    17'b00011011000111101,
    17'b00011011010001111,
    17'b00011011110000101,
    17'b00011100011001101,
    17'b00011110101110001,
    17'b00011110001010010,
    17'b00011100011001101,
    17'b00011101011100001,
    17'b00100010101110001,
    17'b00100101111010111,
    17'b00100111111010111,
    17'b00101000000000000,
    17'b00100111100001010,
    17'b00100100011001101,
    17'b00100000111101100,
    17'b00011101010111000,
    17'b00011010000000000,
    17'b00010101111010111,
    17'b00010010000101001,
    17'b00010000111000011,
    17'b00010000011001101,
    17'b00010011101011100,
    17'b00011000000000000,
    17'b00011110000101001,
    17'b00011011110101110,
    17'b00010111000010100,
    17'b00010101110101110,
    17'b00010110111000011,
    17'b00010111110000101,
    17'b00010111110101110,
    17'b00010111001100110,
    17'b00010111010111000,
    17'b00010111101011100,
    17'b00010111111010111,
    17'b00011000000101001,
    17'b00011000000000000,
    17'b00010110100011111,
    17'b00010100011110110,
    17'b00010010001111011,
    17'b00001111111010111,
    17'b00001101110000101,
    17'b00001100001111011,
    17'b00001011010001111,
    17'b00001011001100110,
    17'b00001011110101110,
    17'b00001100000101001,
    17'b00001101000010100,
    17'b00001101100110011,
    17'b00001101000111101,
    17'b00010100000000000,
    17'b00010110111000011,
    17'b00010010111000011,
    17'b00001110010100100,
    17'b00000110101001000,
    17'b00000010110011010,
    17'b00000000111000011,
    17'b00000000101110001,
    17'b00000001101011100,
    17'b00000011001100110,
    17'b00000011101011100,
    17'b00000010001111011,
    17'b11111111011100001,
    17'b11111110000101001,
    17'b11111100111000011,
    17'b11111011100110011,
    17'b11111011010111000,
    17'b11111011111010111,
    17'b11111101011100001,
    17'b11111111001100110,
    17'b00000101110101110,
    17'b00011000110011010,
    17'b00000000010100100,
    17'b11110111001100110,
    17'b11111011000010100,
    17'b11111100111000011,
    17'b11111011101011100,
    17'b11111011110101110,
    17'b11111011010001111,
    17'b11111100000000000,
    17'b11111011110101110,
    17'b11111010100011111,
    17'b11111000111101100,
    17'b11111001000010100,
    17'b11111101110000101,
    17'b00000001001100110,
    17'b00000011011100001,
    17'b00000100010100100,
    17'b00000100011110110,
    17'b00000011010111000,
    17'b00000000001111011,
    17'b11111101110101110,
    17'b00000000111101100,
    17'b00000100010100100,
    17'b00000110010100100,
    17'b00000110011001101,
    17'b00000101001100110,
    17'b00000011100001010,
    17'b00000001110101110,
    17'b00000010001111011,
    17'b00000001010001111,
    17'b00000010101110001,
    17'b00000100011001101,
    17'b00000010111000011,
    17'b00000001100110011,
    17'b00000011100001010,
    17'b00001000111101100,
    17'b00001101010001111,
    17'b00001101100110011,
    17'b00001011010001111,
    17'b00000111010001111,
    17'b00000101100110011,
    17'b00000101101011100,
    17'b00001000001111011,
    17'b00001101100110011,
    17'b00010010001010010,
    17'b00010101101011100,
    17'b00011000011110110,
    17'b00011100000101001,
    17'b00011100111101100,
    17'b00011100100011111,
    17'b00100000001010010,
    17'b00100001011100001,
    17'b00100010010100100,
    17'b00100010101001000,
    17'b00100011000010100,
    17'b00100011010001111,
    17'b00100011010001111,
    17'b00100011010111000,
    17'b00100011001100110,
    17'b00100100001010010,
    17'b00100101000010100,
    17'b00100110101001000,
    17'b00100111111010111,
    17'b00101000110011010,
    17'b00101001000010100,
    17'b00101000101110001,
    17'b00101001000010100,
    17'b00101001100110011,
    17'b00101010100011111,
    17'b00101010011110110,
    17'b00101010101110001,
    17'b00101011011100001,
    17'b00101100011001101,
    17'b00101101111010111,
    17'b00101111101011100,
    17'b00110001110101110,
    17'b00110100010100100,
    17'b00110110101001000,
    17'b00110110110011010,
    17'b00110111010001111,
    17'b00110111001100110,
    17'b00111000010100100,
    17'b00111000111101100,
    17'b00111001100001010,
    17'b00111011001100110,
    17'b00111101010111000,
    17'b00111101101011100,
    17'b00111101101011100,
    17'b00111101110101110,
    17'b00111101001100110,
    17'b00111101001100110,
    17'b00111101101011100,
    17'b00111110110011010,
    17'b01000000000000000,
    17'b01000000101110001,
    17'b01000001000010100,
    17'b01000001100001010,
    17'b01000010001010010,
    17'b01000010100011111,
    17'b01000010111101100,
    17'b01000010011001101,
    17'b01000001101011100,
    17'b01000000011110110,
    17'b01000000000000000,
    17'b01000000000101001,
    17'b01000001000010100,
    17'b01000010100011111,
    17'b01000100100011111,
    17'b01000110001111011,
    17'b01001000000000000,
    17'b01001010101110001,
    17'b01001101010111000,
    17'b01001110111101100,
    17'b01010001001100110,
    17'b01010010110011010,
    17'b01010011110101110,
    17'b01001100100011111,
    17'b01001011000111101,
    17'b01001010000101001,
    17'b01001010000000000,
    17'b01001010011001101,
    17'b01001010011110110,
    17'b01001010010100100,
    17'b01001010000101001,
    17'b01001001010111000,
    17'b01001001100001010,
    17'b01001010110011010,
    17'b01001100010100100,
    17'b01001110001010010,
    17'b01010000111000011,
    17'b01010010101110001,
    17'b01010100100011111,
    17'b01010110001111011,
    17'b01010111101011100,
    17'b01011000000000000,
    17'b01010111100001010,
    17'b01010111010001111,
    17'b01010110111101100,
    17'b01010110111000011,
    17'b01010110101001000,
    17'b01010110010100100,
    17'b01010110000101001,
    17'b01010101100110011,
    17'b01010101100001010,
    17'b01010101000111101,
    17'b01010101000010100,
    17'b01010100010100100,
    17'b01010011100110011,
    17'b01010010111101100,
    17'b01010011001100110,
    17'b01010100000101001,
    17'b01010100011110110,
    17'b01010100111000011,
    17'b01010100101110001,
    17'b01010011110101110,
    17'b01010010111101100,
    17'b01010010110011010,
    17'b01010010111101100,
    17'b01010011000111101,
    17'b01010011010111000,
    17'b01010011011100001,
    17'b01010011101011100,
    17'b01010011010001111,
    17'b01010011000010100,
    17'b01010010101001000,
    17'b01010010010100100,
    17'b01010001110101110,
    17'b01010001010111000,
    17'b01010000110011010,
    17'b01001110001010010,
    17'b01001101100110011,
    17'b01001101100001010,
    17'b01001101011100001,
    17'b01001101010111000,
    17'b01001100110011010,
    17'b01001100001010010,
    17'b01001011100001010,
    17'b01001010100011111,
    17'b01001001100001010,
    17'b01001000101110001,
    17'b01001000001111011,
    17'b01001000000000000,
    17'b01001000001111011,
    17'b01001000001010010,
    17'b01001000011001101,
    17'b01001000101110001,
    17'b01001001000010100,
    17'b01001001010111000,
    17'b01001001100110011,
    17'b01001001000010100,
    17'b01001000001111011,
    17'b01000111100110011,
    17'b01000101101011100,
    17'b01000011110101110,
    17'b01000011000010100,
    17'b01000011010111000,
    17'b01000110011001101,
    17'b01001000111000011,
    17'b01001011000111101,
    17'b01001100011110110,
    17'b01001101111010111,
    17'b01001111011100001,
    17'b01010000101110001,
    17'b01010001000010100,
    17'b01010000110011010,
    17'b01010001001100110,
    17'b01010001010111000,
    17'b01010001101011100,
    17'b01010000010100100,
    17'b01010010111101100,
    17'b01010100001010010,
    17'b01010011000111101,
    17'b01010001111010111,
    17'b01010001010001111,
    17'b01010001010111000,
    17'b01010001011100001,
    17'b01010001111010111,
    17'b01010001010111000,
    17'b01010100001010010,
    17'b01010111010001111,
    17'b01011001110101110,
    17'b01010110100011111,
    17'b01011101010111000,
    17'b01011100111000011,
    17'b01011010000101001,
    17'b01011111100001010,
    17'b01100011111010111,
    17'b01101100000000000,
    17'b01011000000000000,
    17'b01001001101011100,
    17'b00111111010111000,
    17'b00111000011001101,
    17'b00110010100011111,
    17'b00101110000000000,
    17'b00101101111010111,
    17'b00110000011110110,
    17'b00110110001111011,
    17'b00111100110011010,
    17'b01000100100011111,
    17'b01001000101110001,
    17'b01001011010111000,
    17'b01001110100011111,
    17'b01010000101001000,
    17'b01010001000111101,
    17'b01010000111000011,
    17'b01010001001100110,
    17'b01010010001010010,
    17'b01010011110101110,
    17'b01010100111000011,
    17'b01010101010111000,
    17'b01010101110000101,
    17'b01010101100110011,
    17'b01001001110000101,
    17'b00110011111010111,
    17'b00101000011001101,
    17'b00111000000101001,
    17'b01000001100001010,
    17'b01001001101011100,
    17'b01001101100001010,
    17'b01010001010001111,
    17'b01010100101001000,
    17'b01011000001010010,
    17'b01011001011100001,
    17'b01011001110000101,
    17'b01011000011001101,
    17'b01010011011100001,
    17'b01001001000111101,
    17'b01001001110101110,
    17'b01010011011100001,
    17'b01010011101011100,
    17'b01010010101001000,
    17'b01010001010111000,
    17'b01010000001010010,
    17'b01001110011001101,
    17'b01001100100011111,
    17'b01000011111010111,
    17'b01000001001100110,
    17'b00111011011100001,
    17'b00101111100001010,
    17'b00101111000111101,
    17'b00111010011001101,
    17'b01000110001010010,
    17'b01000101100110011,
    17'b01000011010111000,
    17'b01000011101011100,
    17'b01000010111101100,
    17'b01000011100001010,
    17'b01000101110000101,
    17'b01001111100110011,
    17'b01010010011110110,
    17'b01010000101001000,
    17'b01001101110101110,
    17'b01010011000010100,
    17'b01001100011001101,
    17'b01000011110000101,
    17'b00111111000010100,
    17'b00111111000010100,
    17'b00111101000111101,
    17'b00111111011100001,
    17'b01000110011001101,
    17'b01001100000101001,
    17'b01010010110011010,
    17'b01001111110000101,
    17'b01001011111010111,
    17'b01000101101011100,
    17'b01000001010111000,
    17'b00111101101011100,
    17'b00111010010100100,
    17'b00111000111101100,
    17'b00111000011001101,
    17'b00111000100011111,
    17'b00111000111000011,
    17'b00111001010111000,
    17'b00111001100110011,
    17'b00111010001010010,
    17'b00111011000010100,
    17'b00111010111101100,
    17'b00111010001111011,
    17'b00111001011100001,
    17'b00111000010100100,
    17'b00110111011100001,
    17'b00110110100011111,
    17'b00110101001100110,
    17'b00110100000000000,
    17'b00110011010001111,
    17'b00110011000010100,
    17'b00110011000111101,
    17'b00110100000101001,
    17'b00110100111101100,
    17'b00110110111000011,
    17'b00110111001100110,
    17'b00110110111101100,
    17'b00110110110011010,
    17'b00110110001010010,
    17'b00110101011100001,
    17'b00110100110011010,
    17'b00110100011110110,
    17'b00110011101011100,
    17'b00110011000010100,
    17'b00110010011001101,
    17'b00110010111101100,
    17'b00110011000111101,
    17'b00110010101110001,
    17'b00110010101110001,
    17'b00110010011110110,
    17'b00110010100011111,
    17'b00110010000101001,
    17'b00110001110000101,
    17'b00110000011001101,
    17'b00110000000000000,
    17'b00110000101001000,
    17'b00110000001010010,
    17'b00101110111000011,
    17'b00101101000111101,
    17'b00101011110101110,
    17'b00101010011110110,
    17'b00101001001100110,
    17'b00100111100001010,
    17'b00100101111010111,
    17'b00100100110011010,
    17'b00100011010111000,
    17'b00100011000111101,
    17'b00100011111010111,
    17'b00100101001100110,
    17'b00100110011110110,
    17'b00101011110101110,
    17'b00101100111101100,
    17'b00101001001100110,
    17'b00100100010100100,
    17'b00101000011001101,
    17'b00101011000111101,
    17'b00101100111101100,
    17'b00110001010111000,
    17'b00111010010100100,
    17'b00111010110011010,
    17'b00110110010100100,
    17'b00101111111010111,
    17'b00101110000101001,
    17'b00101000001010010,
    17'b00100000000101001,
    17'b00011110111101100,
    17'b00100010101001000,
    17'b00100010100011111,
    17'b00100101010001111,
    17'b00100011101011100,
    17'b00011110111101100,
    17'b00011101001100110,
    17'b00011111010111000,
    17'b00100001001100110,
    17'b00100001110101110,
    17'b00100100101001000,
    17'b00101000110011010,
    17'b00110000110011010,
    17'b00110011110101110,
    17'b00110100000000000,
    17'b00110010111101100,
    17'b00110010001010010,
    17'b00110000111000011,
    17'b00101111001100110,
    17'b00101011100001010,
    17'b00100111101011100,
    17'b00101001111010111,
    17'b00101011001100110,
    17'b00101100001010010,
    17'b00101110101110001,
    17'b00101111100110011,
    17'b00110010001111011,
    17'b00110010001111011,
    17'b00110100111101100,
    17'b00111001101011100,
    17'b00111011011100001,
    17'b00111011111010111,
    17'b00110111110101110,
    17'b00110110100011111,
    17'b00111001000111101,
    17'b00111100001010010,
    17'b00111000010100100,
    17'b00101111110101110,
    17'b00110001000111101,
    17'b00110101110000101,
    17'b00111000011001101,
    17'b00110110001111011,
    17'b00110110011001101,
    17'b00110100101110001,
    17'b00110111010001111,
    17'b00110110101110001,
    17'b00101111100001010,
    17'b00101011100001010,
    17'b00101111000010100,
    17'b00110010111000011,
    17'b00110101100110011,
    17'b00110100110011010,
    17'b00110110001111011,
    17'b00111001100110011,
    17'b00111110110011010,
    17'b00111011010111000,
    17'b01000110111000011,
    17'b01000111011100001,
    17'b01000110110011010,
    17'b01000100011110110,
    17'b01000110110011010,
    17'b01000101001100110,
    17'b00111111001100110,
    17'b01010010001111011,
    17'b01010010010100100,
    17'b01000001010111000,
    17'b00111000011110110,
    17'b00101111110101110,
    17'b00100100101001000,
    17'b00011000010100100,
    17'b00010010101001000,
    17'b00010101100001010,
    17'b00101000001010010,
    17'b00110101010001111,
    17'b00101101101011100,
    17'b00110001010111000,
    17'b00111100100011111,
    17'b00111110001111011,
    17'b00111001100001010,
    17'b00111000011001101,
    17'b00111010000101001,
    17'b00111101000010100,
    17'b01000101010001111,
    17'b01001001100110011,
    17'b01001101010001111,
    17'b01001101110101110,
    17'b01001011010111000,
    17'b01000101100110011,
    17'b01000001101011100,
    17'b00111110010100100,
    17'b00111001011100001,
    17'b00110101011100001,
    17'b00110100000101001,
    17'b00110100101001000,
    17'b00110110110011010,
    17'b00111001110101110,
    17'b00111010011110110,
    17'b00111011100001010,
    17'b00111100101001000,
    17'b00111100101110001,
    17'b00111011000111101,
    17'b00110110000101001,
    17'b00110111010111000,
    17'b00111001000111101,
    17'b00111011000111101,
    17'b00111100010100100,
    17'b00111101010001111,
    17'b00111100111000011,
    17'b00111101000010100,
    17'b00111110000000000,
    17'b00111111010111000,
    17'b01000000001111011,
    17'b01000000010100100,
    17'b01000001011100001,
    17'b01000001010111000,
    17'b01000000001010010,
    17'b00111110011110110,
    17'b00111100101110001,
    17'b00111010101110001,
    17'b00111010001010010,
    17'b00111000011110110,
    17'b00110110011001101,
    17'b00110110100011111,
    17'b00111001111010111,
    17'b00111110000000000,
    17'b00111111000111101,
    17'b00111110110011010,
    17'b00111101011100001,
    17'b00111110011110110,
    17'b00111110000000000,
    17'b00111101001100110,
    17'b00111000011110110,
    17'b00110111110000101,
    17'b00111010000101001,
    17'b00111011111010111,
    17'b00111011100001010,
    17'b00111001000111101,
    17'b00110110001010010,
    17'b00110011100001010,
    17'b00110001111010111,
    17'b00110000000101001,
    17'b00101110111000011,
    17'b00101110011110110,
    17'b00110010101001000,
    17'b00101110111101100,
    17'b00101101110101110,
    17'b00101111000111101,
    17'b00101111100110011,
    17'b00101110111000011,
    17'b00101110000101001,
    17'b00101101000010100,
    17'b00101101000111101,
    17'b00101010111000011,
    17'b00101001010001111,
    17'b00100111111010111,
    17'b00100111010111000,
    17'b00100111010111000,
    17'b00101010011110110,
    17'b00100111100001010,
    17'b00100110011110110,
    17'b00100110001111011,
    17'b00100100001010010,
    17'b00100010110011010,
    17'b00100011100001010,
    17'b00100000000101001,
    17'b00011100111000011,
    17'b00011100101110001,
    17'b00011111010111000,
    17'b00100011001100110,
    17'b00100100110011010,
    17'b00100011010001111,
    17'b00100001001100110,
    17'b00011111001100110,
    17'b00011101110101110,
    17'b00011101011100001,
    17'b00011110000101001,
    17'b00011110011001101,
    17'b00011101101011100,
    17'b00011100000000000,
    17'b00011001011100001,
    17'b00010111101011100,
    17'b00010110011001101,
    17'b00010101100110011,
    17'b00010101010001111,
    17'b00010100101001000,
    17'b00010010001010010,
    17'b00001111110000101,
    17'b00001101000111101,
    17'b00001000011001101,
    17'b00000101110000101,
    17'b00000010001010010,
    17'b11111110011001101,
    17'b11111011110000101,
    17'b11111000011110110,
    17'b11110111000010100,
    17'b11111010000101001,
    17'b11110111100001010,
    17'b11111001001100110,
    17'b11111100111101100,
    17'b00000010001010010,
    17'b00000101010001111,
    17'b00001000000000000,
    17'b00001011010111000,
    17'b00001100011001101,
    17'b00001100111101100,
    17'b00001100001010010,
    17'b00001001011100001,
    17'b00000111111010111,
    17'b00000101101011100,
    17'b00000111110101110,
    17'b00001000111101100,
    17'b00000111011100001,
    17'b00000110001111011,
    17'b00000110000101001,
    17'b00000101111010111,
    17'b00000100001111011,
    17'b00000000111000011,
    17'b11111111100001010,
    17'b11111101110101110,
    17'b11111101100110011,
    17'b11111101010111000,
    17'b11111101100110011,
    17'b11111100001010010,
    17'b11111001010111000,
    17'b11111001101011100,
    17'b11111010001111011,
    17'b11111011101011100,
    17'b11111100110011010,
    17'b11111111100110011,
    17'b00000100001111011,
    17'b11111111111010111,
    17'b11111111110101110,
    17'b11111111010001111,
    17'b11111101100110011,
    17'b11111100101110001,
    17'b11111000010100100,
    17'b11110010101110001,
    17'b11101111000111101,
    17'b11101111000111101,
    17'b11110000010100100,
    17'b11110100111101100,
    17'b11110100111101100,
    17'b11110110110011010,
    17'b11110111010111000,
    17'b11110111011100001,
    17'b11111000111101100,
    17'b11111011110101110,
    17'b11111101000111101,
    17'b11111100001010010,
    17'b11111111010111000,
    17'b11111101110000101,
    17'b11111010001010010,
    17'b11110110001010010,
    17'b11110001010111000,
    17'b11101011010001111,
    17'b11100100111000011,
    17'b11011110011001101,
    17'b11011000101110001,
    17'b11010100001111011,
    17'b11010100011110110,
    17'b11010011100110011,
    17'b11010101000111101,
    17'b11010110110011010,
    17'b11010110011110110,
    17'b11010111111010111,
    17'b11011001110000101,
    17'b11011010010100100,
    17'b11011011110101110,
    17'b11011101000111101,
    17'b11011110011110110,
    17'b11100000011001101,
    17'b11100010101110001,
    17'b11100100001010010,
    17'b11100100111101100,
    17'b11100101010001111,
    17'b11100101000010100,
    17'b11100100111101100,
    17'b11100101011100001,
    17'b11100110000000000,
    17'b11100110101110001,
    17'b11101000001111011,
    17'b11101010010100100,
    17'b11101100011110110,
    17'b11101110101110001,
    17'b11110000101001000,
    17'b11110011010001111,
    17'b11110001100110011,
    17'b11110101000010100,
    17'b11110011111010111,
    17'b11110100111000011,
    17'b11110101100001010,
    17'b11110101100110011,
    17'b11110101000111101,
    17'b11110101001100110,
    17'b11110101000010100,
    17'b11110100000000000,
    17'b11110011111010111,
    17'b11110101000010100,
    17'b11110010100011111,
    17'b11110100000101001,
    17'b11111101010001111,
    17'b11111110001111011,
    17'b11111101110000101,
    17'b11111100011001101,
    17'b11110001000111101,
    17'b11010011100110011,
    17'b10110111100110011,
    17'b10101001000111101,
    17'b10110000101001000,
    17'b11001111101011100,
    17'b11110101000010100,
    17'b11111011101011100,
    17'b00000011110101110,
    17'b00010000001111011,
    17'b00010111010111000,
    17'b00001111010111000,
    17'b00000011000111101,
    17'b11111011100001010,
    17'b11111000011001101,
    17'b11110100110011010,
    17'b11101101101011100,
    17'b11101001000010100,
    17'b11100110110011010,
    17'b11100110111101100,
    17'b11101000110011010,
    17'b11101010001010010,
    17'b11101011010111000,
    17'b11101011110101110,
    17'b11101011110101110,
    17'b11101010111000011,
    17'b11101001010001111,
    17'b11100111100110011,
    17'b11101000011001101,
    17'b11101010001010010,
    17'b11101010001010010,
    17'b11101000000000000,
    17'b11100111100110011,
    17'b11100100100011111,
    17'b11101000011001101,
    17'b11100110001111011,
    17'b11101001100001010,
    17'b11101010100011111,
    17'b11101100011001101,
    17'b11101001110101110,
    17'b11101001000111101,
    17'b11101001000010100,
    17'b11101011001100110,
    17'b11101100010100100,
    17'b11101010000000000,
    17'b11101111100110011,
    17'b11110011110000101,
    17'b11110100110011010,
    17'b11110101100001010,
    17'b11110101101011100,
    17'b11111000000101001,
    17'b11111010111000011,
    17'b11111100000000000,
    17'b11111100101001000,
    17'b11111101010001111,
    17'b11111101110101110,
    17'b11111110011001101,
    17'b11111110011001101,
    17'b11111101111010111,
    17'b11111100010100100,
    17'b11111010011001101,
    17'b11111000010100100,
    17'b11110110010100100,
    17'b11110100000101001,
    17'b11110010100011111,
    17'b11110001111010111,
    17'b11110001010111000,
    17'b11110001110000101,
    17'b11110010011001101,
    17'b11110011001100110,
    17'b11110100001010010,
    17'b11110101100001010,
    17'b11111000011110110,
    17'b11111010111000011,
    17'b11111101100001010,
    17'b11111110110011010,
    17'b11111111011100001,
    17'b11111111001100110,
    17'b11111110100011111,
    17'b11111101011100001,
    17'b11111011101011100,
    17'b11111001100001010,
    17'b11111000000101001,
    17'b11110110110011010,
    17'b11110101110101110,
    17'b11110100110011010,
    17'b11110011011100001,
    17'b11110010001111011,
    17'b11110000101110001,
    17'b11101111011100001,
    17'b11101110011001101,
    17'b11101110011001101,
    17'b11101110001010010,
    17'b11101101100001010,
    17'b11101101001100110,
    17'b11101101101011100,
    17'b11101110111000011,
    17'b11110000101110001,
    17'b11110000101001000,
    17'b11110000001111011,
    17'b11101111101011100,
    17'b11110000010100100,
    17'b11110000001111011,
    17'b11110000111101100,
    17'b11110001101011100,
    17'b11110010001111011,
    17'b11110100010100100,
    17'b11110100011001101,
    17'b11110011101011100,
    17'b11110010101110001,
    17'b11110001110000101,
    17'b11101110010100100,
    17'b11101101110101110,
    17'b11101101110000101,
    17'b11101100001111011,
    17'b11101011010111000,
    17'b11101011011100001,
    17'b11101011101011100,
    17'b11101011001100110,
    17'b11101010101110001,
    17'b11101010000101001,
    17'b11101001100110011,
    17'b11101001010001111,
    17'b11101001000111101,
    17'b11101001010001111,
    17'b11101001011100001,
    17'b11101001110000101,
    17'b11101001110000101,
    17'b11101010000000000,
    17'b11101010000101001,
    17'b11101010011110110,
    17'b11101010101110001,
    17'b11101011000111101,
    17'b11101011010001111,
    17'b11101011001100110,
    17'b11101011010111000,
    17'b11101011011100001,
    17'b11101011100110011,
    17'b11101011100110011,
    17'b11101011110101110,
    17'b11101100001010010,
    17'b11101100100011111,
    17'b11101100101001000,
    17'b11101100011110110,
    17'b11101100001111011,
    17'b11101100000000000,
    17'b11101011010001111,
    17'b11101010000101001,
    17'b11101001010111000,
    17'b11101000101001000,
    17'b11101000010100100,
    17'b11101000011110110,
    17'b11101001010111000,
    17'b11101001110000101,
    17'b11101001110000101,
    17'b11101001110000101,
    17'b11101001100001010,
    17'b11101010000000000,
    17'b11101010110011010,
    17'b11101011100110011,
    17'b11101100000101001,
    17'b11101101100110011,
    17'b11110100000000000,
    17'b11110100101110001,
    17'b11110011011100001,
    17'b11110001001100110,
    17'b11101101101011100,
    17'b11101010101110001,
    17'b11101001010001111,
    17'b11101010000101001,
    17'b11101011111010111,
    17'b11101101100001010,
    17'b11101110011001101,
    17'b11101110000101001,
    17'b11101101010111000,
    17'b11101101010111000,
    17'b11101101101011100,
    17'b11101110111101100,
    17'b11101111110101110,
    17'b11110000000101001,
    17'b11101111110101110,
    17'b11101111101011100,
    17'b11101111010001111,
    17'b11101110000101001,
    17'b11101101000111101,
    17'b11101100101110001,
    17'b11101100010100100,
    17'b11101011101011100,
    17'b11101010001010010,
    17'b11101000111101100,
    17'b11100111010111000,
    17'b11100110011001101,
    17'b11100101100110011,
    17'b11100101000111101,
    17'b11100100111101100,
    17'b11100011000111101,
    17'b11100011111010111,
    17'b11100100011001101,
    17'b11100100001111011,
    17'b11100011111010111,
    17'b11100011001100110,
    17'b11100010010100100,
    17'b11100000011110110,
    17'b11011110011001101,
    17'b11011010010100100,
    17'b11011011010001111,
    17'b11011011000010100,
    17'b11011011001100110,
    17'b11011010110011010,
    17'b11011010011110110,
    17'b11011011110000101,
    17'b11011100011110110,
    17'b11011110000101001,
    17'b11011111011100001,
    17'b11100000110011010,
    17'b11100001010111000,
    17'b11100010010100100,
    17'b11100011010001111,
    17'b11100101001100110,
    17'b11100111011100001,
    17'b11101001010001111,
    17'b11101011000111101,
    17'b11101101010111000,
    17'b11101110101110001,
    17'b11110000000000000,
    17'b11110000101110001,
    17'b11110001010001111,
    17'b11110001100110011,
    17'b11110010010100100,
    17'b11110010010100100,
    17'b11110010000000000,
    17'b11110001011100001,
    17'b11110000111000011,
    17'b11110000010100100,
    17'b11101110110011010,
    17'b11101100101110001,
    17'b11101011000010100,
    17'b11100101110000101,
    17'b11011010011110110,
    17'b11100000010100100,
    17'b11100101110101110,
    17'b11101001100110011,
    17'b11110000101001000,
    17'b11111000010100100,
    17'b11111111111010111,
    17'b00000111011100001,
    17'b00000110111101100,
    17'b00000010011110110,
    17'b00000011000010100,
    17'b00000010000101001,
    17'b00000010111000011,
    17'b00000001000111101,
    17'b00000010010100100,
    17'b00000001110101110,
    17'b00000000001010010,
    17'b00000001011100001,
    17'b00000100000000000,
    17'b00000101001100110,
    17'b00000101110101110,
    17'b00000101010001111,
    17'b00000111010001111,
    17'b00001100011110110,
    17'b00001101110000101,
    17'b00010000100011111,
    17'b00010011001100110,
    17'b00010101110000101,
    17'b00010111011100001,
    17'b00011000010100100,
    17'b00011000011001101,
    17'b00011000101001000,
    17'b00011000010100100,
    17'b00010111010111000,
    17'b00010110010100100,
    17'b00010101000111101,
    17'b00010011100110011,
    17'b00010010101110001,
    17'b00010010001010010,
    17'b00010001010001111,
    17'b00010000100011111,
    17'b00010000100011111,
    17'b00010001101011100,
    17'b00010011000111101,
    17'b00010011111010111,
    17'b00010101100110011,
    17'b00010111010111000,
    17'b00010111001100110,
    17'b00010100011110110,
    17'b00010001101011100,
    17'b00010000000101001,
    17'b00010000011110110,
    17'b00010001010111000,
    17'b00010010001111011,
    17'b00010010011110110,
    17'b00010010100011111,
    17'b00010010010100100,
    17'b00010001101011100,
    17'b00010001010111000,
    17'b00010001000111101,
    17'b00010001010001111,
    17'b00010001000111101,
    17'b00010001001100110,
    17'b00010001100110011,
    17'b00010001011100001,
    17'b00010000111101100,
    17'b00010000101110001,
    17'b00010000011001101,
    17'b00010000110011010,
    17'b00010001010111000,
    17'b00010011010001111,
    17'b00010011111010111,
    17'b00010010011001101,
    17'b00010000111101100,
    17'b00010000000101001,
    17'b00001111010111000,
    17'b00001110100011111,
    17'b00001101110101110,
    17'b00001101101011100,
    17'b00001110101001000,
    17'b00001111011100001,
    17'b00010000000101001,
    17'b00010000011110110,
    17'b00010000011001101,
    17'b00001111110101110,
    17'b00001110100011111,
    17'b00001101000010100,
    17'b00001011110101110,
    17'b00001011000010100,
    17'b00001010011001101,
    17'b00001001100110011,
    17'b00001000111101100,
    17'b00001000100011111,
    17'b00000111111010111,
    17'b00000110011001101,
    17'b11111111100001010,
    17'b11111110001010010,
    17'b11111100101001000,
    17'b11111011100001010,
    17'b11111010001010010,
    17'b11111001010001111,
    17'b11111000110011010,
    17'b11110110011110110,
    17'b11111111100110011,
    17'b00001011101011100,
    17'b00001100000000000,
    17'b00001001110101110,
    17'b00000011010111000,
    17'b11111011010111000,
    17'b11111000001010010,
    17'b11110101100110011,
    17'b11110010011110110,
    17'b11110001110101110,
    17'b11110001001100110,
    17'b11101101010111000,
    17'b11101100000000000,
    17'b11101011000111101,
    17'b11100101100001010,
    17'b11100100111101100,
    17'b11101100001111011,
    17'b11110000110011010,
    17'b11110010000000000,
    17'b11110010000000000,
    17'b11110010101001000,
    17'b11110100000101001,
    17'b11110110101110001,
    17'b11111010001111011,
    17'b11111110111000011,
    17'b00000010111000011,
    17'b00001000000101001,
    17'b00000110010100100,
    17'b00000100000101001,
    17'b00000001000111101,
    17'b11111100000000000,
    17'b11111000011110110,
    17'b11110110000000000,
    17'b11110100000000000,
    17'b11110010000101001,
    17'b11110000110011010,
    17'b11101111111010111,
    17'b11101111101011100,
    17'b11101111111010111,
    17'b11110000010100100,
    17'b11110000001111011,
    17'b11110000011110110,
    17'b11110010001111011,
    17'b11110011111010111,
    17'b11110100111101100,
    17'b11110101011100001,
    17'b11110101000111101,
    17'b11110100101001000,
    17'b11110100000101001,
    17'b11110011011100001,
    17'b11110011100001010,
    17'b11110011110101110,
    17'b11110100101001000,
    17'b11110101110101110,
    17'b11110111001100110,
    17'b11111000001010010,
    17'b11111001100001010,
    17'b11111011110000101,
    17'b11111100111000011,
    17'b11111110110011010,
    17'b00000000111000011,
    17'b00000010111000011,
    17'b00000100000000000,
    17'b00000101010001111,
    17'b00000110111000011,
    17'b00001000001010010,
    17'b00001000001010010,
    17'b00000111100001010,
    17'b00000111110000101,
    17'b00001000000000000,
    17'b00001000111000011,
    17'b00001001110101110,
    17'b00001010110011010,
    17'b00001010001111011,
    17'b00001001100110011,
    17'b00001000100011111,
    17'b00000111000010100,
    17'b00000101011100001,
    17'b00000011101011100,
    17'b00000011010111000,
    17'b00000010000101001,
    17'b00000000000000000,
    17'b11111110001010010,
    17'b11111101000010100,
    17'b11111011001100110,
    17'b11111010010100100,
    17'b11111100001111011,
    17'b11111101111010111,
    17'b11111110010100100,
    17'b11111101101011100,
    17'b11111100111000011,
    17'b11111101010001111,
    17'b11111110001111011,
    17'b11111111101011100,
    17'b00000001110101110,
    17'b00000011000010100,
    17'b00000100010100100,
    17'b00000101110101110,
    17'b00000110101001000,
    17'b00000111011100001,
    17'b00000111111010111,
    17'b00000111010001111,
    17'b00000110010100100,
    17'b00000101000111101,
    17'b00000100000000000,
    17'b00000011111010111,
    17'b00000011110101110,
    17'b00000011100110011,
    17'b00000100010100100,
    17'b00000101001100110,
    17'b00000101000111101,
    17'b00000100101110001,
    17'b00000011011100001,
    17'b00000000101110001,
    17'b11111110011001101,
    17'b11111101001100110,
    17'b11111100101110001,
    17'b11111100010100100,
    17'b11111100001111011,
    17'b11111101010001111,
    17'b11111111010001111,
    17'b00000001000010100,
    17'b00000010111000011,
    17'b00000011011100001,
    17'b00000011101011100,
    17'b00000011010111000,
    17'b00000010000000000,
    17'b00000000011110110,
    17'b11111111100001010,
    17'b11111110110011010,
    17'b11111101101011100,
    17'b11111101001100110,
    17'b11111100010100100,
    17'b11111010010100100,
    17'b11111001100001010,
    17'b11111001111010111,
    17'b11110101010001111,
    17'b11111001010111000,
    17'b11111100001111011,
    17'b11111101000010100,
    17'b11111101001100110,
    17'b11111101101011100,
    17'b11110011100001010,
    17'b11111000101110001,
    17'b11111110101001000,
    17'b11111101111010111,
    17'b11111100001010010,
    17'b11111010111000011,
    17'b11110111000111101,
    17'b11110101000111101,
    17'b11110101111010111,
    17'b11110110000000000,
    17'b11110101101011100,
    17'b11110101100110011,
    17'b11110101000010100,
    17'b11110100101001000,
    17'b11110101000010100,
    17'b11110110001111011,
    17'b11110110111000011,
    17'b11111000000000000,
    17'b11111000000000000,
    17'b11110110101001000,
    17'b11110101110101110,
    17'b11110011111010111,
    17'b11110011111010111,
    17'b11110100101001000,
    17'b11110010000101001,
    17'b11101111100110011,
    17'b11110000010100100,
    17'b11110010111000011,
    17'b11110001011100001,
    17'b11110011010111000,
    17'b11110001101011100,
    17'b11101110110011010,
    17'b11101010001111011,
    17'b11101101100110011,
    17'b11110011010111000,
    17'b11110101000010100,
    17'b11110111110000101,
    17'b11111010000101001,
    17'b11110111110101110,
    17'b11110101000111101,
    17'b11110011100110011,
    17'b11110010110011010,
    17'b11110000001111011,
    17'b11101110000000000,
    17'b11101100100011111,
    17'b11101011110101110,
    17'b11101011011100001,
    17'b11101001101011100,
    17'b11101001001100110,
    17'b11100110111000011,
    17'b11100111001100110,
    17'b11101000100011111,
    17'b11100111110000101,
    17'b11100110111101100,
    17'b11100110001010010,
    17'b11100101111010111,
    17'b11100101111010111,
    17'b11100110011110110,
    17'b11100110100011111,
    17'b11100110010100100,
    17'b11100101110000101,
    17'b11100110001010010,
    17'b11100111010111000,
    17'b11101000100011111,
    17'b11101001110101110,
    17'b11101010010100100,
    17'b11101011000111101,
    17'b11101011000010100,
    17'b11101010101001000,
    17'b11101010101110001,
    17'b11101001001100110,
    17'b11100111100001010,
    17'b11100101000010100,
    17'b11100011101011100,
    17'b11100001110101110,
    17'b11100000101001000,
    17'b11100000110011010,
    17'b11100010011001101,
    17'b11100001011100001,
    17'b11100000101001000,
    17'b11011111100001010,
    17'b11011111000010100,
    17'b11011110010100100,
    17'b11011110000000000,
    17'b11011101100110011,
    17'b11011100101001000,
    17'b11011011100110011,
    17'b11011011001100110,
    17'b11011011110101110,
    17'b11011011100001010,
    17'b11011010100011111,
    17'b11011010011001101,
    17'b11011010011110110,
    17'b11011100001010010,
    17'b11011100101110001,
    17'b11011101100001010,
    17'b11011111000010100,
    17'b11011111110000101,
    17'b11100001000010100,
    17'b11100001110000101,
    17'b11100001110101110,
    17'b11100001000010100,
    17'b11011111111010111,
    17'b11100000000101001,
    17'b11011111000111101,
    17'b11011101110000101,
    17'b11011100111000011,
    17'b11011101101011100,
    17'b11011110101110001,
    17'b11100000001111011,
    17'b11100000001010010,
    17'b11100000001010010,
    17'b11100010011001101,
    17'b11100100111000011,
    17'b11100111000111101,
    17'b11101011011100001,
    17'b11101110000101001,
    17'b11101111110101110,
    17'b11110001000010100,
    17'b11110010101001000,
    17'b11110011010111000,
    17'b11110100011001101,
    17'b11110100001010010,
    17'b11110100011001101,
    17'b11110100100011111,
    17'b11110011111010111,
    17'b11110010001111011,
    17'b11110000101110001,
    17'b11110000100011111,
    17'b11110001010111000,
    17'b11110010111101100,
    17'b11110100011001101,
    17'b11110101111010111,
    17'b11110111000111101,
    17'b11111000101110001,
    17'b11111001101011100,
    17'b11111010111101100,
    17'b11111100011110110,
    17'b11111110001010010,
    17'b11111111001100110,
    17'b11111111100110011,
    17'b00000000100011111,
    17'b00000001000111101,
    17'b00000001100001010,
    17'b00000001101011100,
    17'b00000001100110011,
    17'b00000000111101100,
    17'b00000000111000011,
    17'b00000001000111101,
    17'b00000001100001010,
    17'b00000010110011010,
    17'b00000011001100110,
    17'b00000011101011100,
    17'b00000100100011111,
    17'b00000101110101110,
    17'b00000111100110011,
    17'b00001000001111011,
    17'b00001000100011111,
    17'b00001000010100100,
    17'b00001000001010010,
    17'b00000111111010111,
    17'b00001000000000000,
    17'b00000111100110011,
    17'b00000110111101100,
    17'b00000110101110001,
    17'b00000110001111011,
    17'b00000101110000101,
    17'b00000101011100001,
    17'b00000101100110011,
    17'b00000101110000101,
    17'b00000101010001111,
    17'b00000100011110110,
    17'b00000011110000101,
    17'b00000000101110001,
    17'b00000000000000000,
    17'b00000010101110001,
    17'b00001000001111011,
    17'b00001110011110110,
    17'b00010000100011111,
    17'b00001110101001000,
    17'b00001100101001000,
    17'b00001100011001101,
    17'b00001100000000000,
    17'b00001101110101110,
    17'b00010000000000000,
    17'b00010001111010111,
    17'b00010011100110011,
    17'b00010100011001101,
    17'b00010100101001000,
    17'b00010100001111011,
    17'b00010100011110110,
    17'b00010100011110110,
    17'b00010100010100100,
    17'b00010011110101110,
    17'b00010011101011100,
    17'b00010011000111101,
    17'b00010010111101100,
    17'b00010011001100110,
    17'b00010011000111101,
    17'b00010011000010100,
    17'b00010010111000011,
    17'b00010011000111101,
    17'b00010011010111000,
    17'b00010011111010111,
    17'b00010100001111011,
    17'b00010100100011111,
    17'b00010100100011111,
    17'b00010011111010111,
    17'b00010011010001111,
    17'b00010010111101100,
    17'b00010010111000011,
    17'b00010010110011010,
    17'b00010011000010100,
    17'b00010011010001111,
    17'b00010011100001010,
    17'b00010011010111000,
    17'b00010011011100001,
    17'b00010010111101100,
    17'b00010010001111011,
    17'b00010001100001010,
    17'b00010000101110001,
    17'b00010001000010100,
    17'b00010001100110011,
    17'b00010010011110110,
    17'b00010011011100001,
    17'b00010011110101110,
    17'b00010100010100100,
    17'b00010100101110001,
    17'b00010101010001111,
    17'b00010100011110110,
    17'b00010100001010010,
    17'b00010011101011100,
    17'b00010000110011010,
    17'b00010000001111011,
    17'b00001111100001010,
    17'b00001111000111101,
    17'b00001111010111000,
    17'b00001111100001010,
    17'b00001111101011100,
    17'b00001111110101110,
    17'b00010000101110001,
    17'b00010001100110011,
    17'b00010010000101001,
    17'b00010010011110110,
    17'b00010010100011111,
    17'b00010011000111101,
    17'b00010011001100110,
    17'b00010011101011100,
    17'b00010011111010111,
    17'b00010011110101110,
    17'b00010011011100001,
    17'b00010010111000011,
    17'b00010010101001000,
    17'b00010010000101001,
    17'b00010010000000000,
    17'b00010001110000101,
    17'b00010001111010111,
    17'b00010010001010010,
    17'b00010010100011111,
    17'b00010010011001101,
    17'b00010001110000101,
    17'b00010001001100110,
    17'b00010000100011111,
    17'b00001111111010111,
    17'b00001111010111000,
    17'b00001111010111000,
    17'b00001111010001111,
    17'b00001111010001111,
    17'b00001111000111101,
    17'b00001110110011010,
    17'b00001110100011111,
    17'b00001110101001000,
    17'b00001111000010100,
    17'b00001111000010100,
    17'b00001111010001111,
    17'b00001111011100001,
    17'b00010000000101001,
    17'b00010000011001101,
    17'b00010000111101100,
    17'b00010001010111000,
    17'b00010001111010111,
    17'b00010010101110001,
    17'b00010011110000101,
    17'b00010011010001111,
    17'b00010010101001000,
    17'b00010001001100110,
    17'b00001110011110110,
    17'b00001011010111000,
    17'b00001010101110001,
    17'b00001010101110001,
    17'b00000101000111101,
    17'b00011101110000101,
    17'b00101001010111000,
    17'b00010110000000000,
    17'b00001101000111101,
    17'b00001010100011111,
    17'b00001001011100001,
    17'b00001001110000101,
    17'b00001001010001111,
    17'b00001001000010100,
    17'b00001010001111011,
    17'b00001011010001111,
    17'b00001100000000000,
    17'b00001011100110011,
    17'b00001010101110001,
    17'b00001001111010111,
    17'b00001001011100001,
    17'b00001001010111000,
    17'b00001001100110011,
    17'b00001010001111011,
    17'b00001010110011010,
    17'b00001010111000011,
    17'b00001010100011111,
    17'b00001010101001000,
    17'b00001010101001000,
    17'b00001010101001000,
    17'b00001010111000011,
    17'b00001010101001000,
    17'b00001001010111000,
    17'b00001001010001111,
    17'b00001001010111000,
    17'b00001001111010111,
    17'b00001010011110110,
    17'b00001010011001101,
    17'b00001010001010010,
    17'b00001010010100100,
    17'b00001010111101100,
    17'b00001011000010100,
    17'b00001011001100110,
    17'b00001010101110001,
    17'b00001010101001000,
    17'b00001010101001000,
    17'b00001010101001000,
    17'b00001001111010111,
    17'b00001001000010100,
    17'b00001000010100100,
    17'b00000110111101100,
    17'b00000101000111101,
    17'b00000011010001111,
    17'b00000001111010111,
    17'b00000001000010100,
    17'b00000000000101001,
    17'b11111111011100001,
    17'b11111110111101100,
    17'b11111111100001010,
    17'b11111111100001010,
    17'b11111111010001111,
    17'b11111110100011111,
    17'b11111101101011100,
    17'b11111100011001101,
    17'b11111011100001010,
    17'b11111011001100110,
    17'b11111011000010100,
    17'b11111011000111101,
    17'b11111011001100110,
    17'b11111011111010111,
    17'b11111100111000011,
    17'b00000100101110001,
    17'b00000111101011100,
    17'b00001100010100100,
    17'b00010000001010010,
    17'b00010100101110001,
    17'b00011000111101100,
    17'b00011110001111011,
    17'b00100001000111101,
    17'b00100010011110110,
    17'b00100010000000000,
    17'b00100000110011010,
    17'b00011110101110001,
    17'b00011100000000000,
    17'b00010111110000101,
    17'b00010100010100100,
    17'b00010001001100110,
    17'b00001101101011100,
    17'b00001010010100100,
    17'b00000110111000011,
    17'b00000101110101110,
    17'b00000100111101100,
    17'b00000100011001101,
    17'b00000100011110110,
    17'b00000100110011010,
    17'b00000100110011010,
    17'b00000100100011111,
    17'b00000100111000011,
    17'b00000100101001000,
    17'b00000100100011111,
    17'b00000101001100110,
    17'b00000110011001101,
    17'b00000111011100001,
    17'b00001000010100100,
    17'b00001001100110011,
    17'b00001010111000011,
    17'b00001100001111011,
    17'b00001101111010111,
    17'b00010000010100100,
    17'b00010001000111101,
    17'b00010001000111101,
    17'b00010000110011010,
    17'b00010000001010010,
    17'b00001111101011100,
    17'b00001111111010111,
    17'b00010000111000011,
    17'b00010000001111011,
    17'b00001111111010111,
    17'b00001111001100110,
    17'b00001110100011111,
    17'b00001100111101100,
    17'b00001011100001010,
    17'b00001010001010010,
    17'b00001001001100110,
    17'b00001000101110001,
    17'b00000111010111000,
    17'b00000101110101110,
    17'b00000100111000011,
    17'b00000100011110110,
    17'b00000100001010010,
    17'b00000101100110011,
    17'b00000110101110001,
    17'b00000111000111101,
    17'b00001000000101001,
    17'b00001000001010010,
    17'b00001000110011010,
    17'b00001001110000101,
    17'b00001010011110110,
    17'b00001011000111101,
    17'b00001011100110011,
    17'b00001011010111000,
    17'b00001100000101001,
    17'b00001011100001010,
    17'b00001001110000101,
    17'b00000111000111101,
    17'b00000101001100110,
    17'b00000011110000101,
    17'b00000010011001101,
    17'b00000010101110001,
    17'b00000001111010111,
    17'b00000000010100100,
    17'b11111110111000011,
    17'b11111111101011100,
    17'b00000000000101001,
    17'b11111111000010100,
    17'b11111110011001101,
    17'b11111101000111101,
    17'b11111100001111011,
    17'b11111100101110001,
    17'b11111101010111000,
    17'b11111110010100100,
    17'b11111111000010100,
    17'b11111111010001111,
    17'b11111111101011100,
    17'b00000001100110011,
    17'b00000101001100110,
    17'b00000011100110011,
    17'b00000010000000000,
    17'b11111101101011100,
    17'b11111100000101001,
    17'b11111001111010111,
    17'b11110110011001101,
    17'b11110110101110001,
    17'b11110110111101100,
    17'b11110101000111101,
    17'b11110010100011111,
    17'b11110000111101100,
    17'b11101111010001111,
    17'b11101111010001111,
    17'b11110000001010010,
    17'b11110001111010111,
    17'b11110011011100001,
    17'b11110100010100100,
    17'b11110100100011111,
    17'b11110011011100001,
    17'b11110010101001000,
    17'b11110001011100001,
    17'b11110000101001000,
    17'b11110000000000000,
    17'b11101111101011100,
    17'b11101111010001111,
    17'b11101111010111000,
    17'b11110000011110110,
    17'b11110001101011100,
    17'b11110011001100110,
    17'b11110100101110001,
    17'b11110110101110001,
    17'b11110111111010111,
    17'b11111000000101001,
    17'b11110110101110001,
    17'b11110100101110001,
    17'b11110010111000011,
    17'b11110001001100110,
    17'b11110000010100100,
    17'b11101111100110011,
    17'b11101110011110110,
    17'b11101101000010100,
    17'b11101011011100001,
    17'b11101010111000011,
    17'b11101010111101100,
    17'b11101011010001111,
    17'b11101010111101100,
    17'b11101010001111011,
    17'b11101001011100001,
    17'b11101001001100110,
    17'b11101001010111000,
    17'b11101010000101001,
    17'b11101010010100100,
    17'b11101110011001101,
    17'b11110100100011111,
    17'b11110000111000011,
    17'b11101010000000000,
    17'b11101111110000101,
    17'b11110011100110011,
    17'b11110101010111000,
    17'b11110100100011111,
    17'b11110011001100110,
    17'b11110011001100110,
    17'b11110100111101100,
    17'b11110110011001101,
    17'b11110111000010100,
    17'b11110110111000011,
    17'b11110101101011100,
    17'b11110010110011010,
    17'b11110000010100100,
    17'b11101101100110011,
    17'b11101011000111101,
    17'b11100111110000101,
    17'b11100110001010010,
    17'b11100101001100110,
    17'b11100100011110110,
    17'b11100011001100110,
    17'b11100010101001000,
    17'b11100010011110110,
    17'b11100010100011111,
    17'b11100010011110110,
    17'b11100001111010111,
    17'b11100001111010111,
    17'b11100001110101110,
    17'b11100001111010111,
    17'b11100010001010010,
    17'b11100011010111000,
    17'b11100100111000011,
    17'b11100110111101100,
    17'b11101000110011010,
    17'b11101001100110011,
    17'b11101010011001101,
    17'b11101011000010100,
    17'b11101011010001111,
    17'b11101010010100100,
    17'b11101001000010100,
    17'b11100111100001010,
    17'b11100101100001010,
    17'b11100100100011111,
    17'b11100011001100110,
    17'b11100001110101110,
    17'b11011111011100001,
    17'b11011101010001111,
    17'b11011010110011010,
    17'b11011000110011010,
    17'b11010111010001111,
    17'b11010100111000011,
    17'b11010011011100001,
    17'b11010010000101001,
    17'b11010000111101100,
    17'b11001111100110011,
    17'b11001111010001111,
    17'b11001111000010100,
    17'b11001110101110001,
    17'b11001110101001000,
    17'b11001110100011111,
    17'b11001110100011111,
    17'b11001110001010010,
    17'b11001101111010111,
    17'b11001101101011100,
    17'b11001101100110011,
    17'b11001101000111101,
    17'b11001100101110001,
    17'b11001100000000000,
    17'b11001010111101100,
    17'b11001010110011010,
    17'b11001010110011010,
    17'b11001011000111101,
    17'b11001011010111000,
    17'b11001011110101110,
    17'b11001011110101110,
    17'b11001010101001000,
    17'b11001001001100110,
    17'b11000111110101110,
    17'b11000011101011100,
    17'b11000010011110110,
    17'b11000001011100001,
    17'b11000000111101100,
    17'b11000000111101100,
    17'b11000001010111000,
    17'b11000010000101001,
    17'b11000010100011111,
    17'b11000011011100001,
    17'b11000100001010010,
    17'b11000101000010100,
    17'b11000101001100110,
    17'b11000101000111101,
    17'b11000100110011010,
    17'b11000011111010111,
    17'b11000010101001000,
    17'b11000000110011010,
    17'b10111111111010111,
    17'b10111111000010100,
    17'b10111110101001000,
    17'b10111110010100100,
    17'b10111110000101001,
    17'b10111101111010111,
    17'b10111101110101110,
    17'b10111110001010010,
    17'b10111110000101001,
    17'b10111101110000101,
    17'b10111101000010100,
    17'b10111100011110110,
    17'b10111011011100001,
    17'b10111010001111011,
    17'b10111000101110001,
    17'b10110111101011100,
    17'b10110110101110001,
    17'b10110101110000101,
    17'b10110101011100001,
    17'b10110101110101110,
    17'b10111000011001101,
    17'b10111001010001111,
    17'b10111001010001111,
    17'b10111001110101110,
    17'b10111010000000000,
    17'b10111100110011010,
    17'b10111101001100110,
    17'b10111101000010100,
    17'b10111101000010100,
    17'b10111101010111000,
    17'b10111101001100110,
    17'b10111101100001010,
    17'b10111101100001010,
    17'b10111100011001101,
    17'b10111011000010100,
    17'b10111010000000000,
    17'b10111001001100110,
    17'b10111001000010100,
    17'b10111001101011100,
    17'b10111010100011111,
    17'b10111011110000101,
    17'b10111100011001101,
    17'b10111101000111101,
    17'b10111101010111000,
    17'b10111101111010111,
    17'b10111110011001101,
    17'b10111111001100110,
    17'b10111111001100110,
    17'b10111110110011010,
    17'b10111110010100100,
    17'b10111101100110011,
    17'b10111100110011010,
    17'b10111100001111011,
    17'b10111100001010010,
    17'b10111100000000000,
    17'b10111100000000000,
    17'b10111011110101110,
    17'b10111100000000000,
    17'b10111100111000011,
    17'b10111101000010100,
    17'b10111101010001111,
    17'b10111101110101110,
    17'b10111110000000000,
    17'b10111110011001101,
    17'b10111111000010100,
    17'b10111111100001010,
    17'b11000000000000000,
    17'b11000000010100100,
    17'b11000000111101100,
    17'b11000001010001111,
    17'b11000010000000000,
    17'b11000010101001000,
    17'b11000011110000101,
    17'b11000100111101100,
    17'b11000101101011100,
    17'b11000110101001000,
    17'b11000111100110011,
    17'b11001000101110001,
    17'b11001001010111000,
    17'b11001010001111011,
    17'b11001011000010100,
    17'b11001011101011100,
    17'b11001100001010010,
    17'b11001100011001101,
    17'b11001100001111011,
    17'b11001011001100110,
    17'b11001010000000000,
    17'b11000111111010111,
    17'b11000110101001000,
    17'b11000000101001000,
    17'b11000000011001101,
    17'b11000000011001101,
    17'b11000000110011010,
    17'b11000001100110011,
    17'b11000010100011111,
    17'b11000011100001010,
    17'b11000100010100100,
    17'b11000101010001111,
    17'b11000101111010111,
    17'b11000110010100100,
    17'b11000110101110001,
    17'b11000111011100001,
    17'b11000111110101110,
    17'b11000111111010111,
    17'b11000111011100001,
    17'b11000111000111101,
    17'b11000110011110110,
    17'b11000101100001010,
    17'b11000100011001101,
    17'b11000011010111000,
    17'b11000010100011111,
    17'b11000000111101100,
    17'b11000000000000000,
    17'b10111110111000011,
    17'b10111110000000000,
    17'b10111101010001111,
    17'b10111100111000011,
    17'b10111100111101100,
    17'b10111100101110001,
    17'b10111101010001111,
    17'b11000101000010100,
    17'b11000101110101110,
    17'b11000101010001111,
    17'b11000101100001010,
    17'b11000110010100100,
    17'b11000111111010111,
    17'b11001000100011111,
    17'b11001001111010111,
    17'b11001010100011111,
    17'b11001100011001101,
    17'b11001101011100001,
    17'b11001111010001111,
    17'b11001110111000011,
    17'b11010000111000011,
    17'b11010010001010010,
    17'b11010010001111011,
    17'b11010011111010111,
    17'b11010100000101001,
    17'b11010100111000011,
    17'b11010101010111000,
    17'b11010110001111011,
    17'b11010110111101100,
    17'b11010111010111000,
    17'b11010111101011100,
    17'b11010111100110011,
    17'b11010111110101110,
    17'b11010111101011100,
    17'b11010111001100110,
    17'b11010110010100100,
    17'b11010101011100001,
    17'b11010100100011111,
    17'b11010100001010010,
    17'b11010100011110110,
    17'b11010101001100110,
    17'b11010110001010010,
    17'b11010111000010100,
    17'b11010111100110011,
    17'b11011000000000000,
    17'b11010111111010111,
    17'b11010111100110011,
    17'b11010111110000101,
    17'b11011000010100100,
    17'b11011001000111101,
    17'b11011010000000000,
    17'b11011011001100110,
    17'b11011100101001000,
    17'b11011101100110011,
    17'b11011110001111011,
    17'b11011110101001000,
    17'b11011110101110001,
    17'b11011101110101110,
    17'b11011100011110110,
    17'b11011010000101001,
    17'b11011000101001000,
    17'b11010110110011010,
    17'b11010100011001101,
    17'b11010010101110001,
    17'b11010001100001010,
    17'b11010000101110001,
    17'b11010000101110001,
    17'b11010001010111000,
    17'b11010100000101001,
    17'b11010101011100001,
    17'b11010111011100001,
    17'b11011001110101110,
    17'b11011011111010111,
    17'b11011101000111101,
    17'b11011101001100110,
    17'b11011101100110011,
    17'b11011100111000011,
    17'b11011111001100110,
    17'b11100010010100100,
    17'b11100100111101100,
    17'b11100111111010111,
    17'b11100111111010111,
    17'b11100110111101100,
    17'b11100101100110011,
    17'b11100101011100001,
    17'b11100101010001111,
    17'b11100100111000011,
    17'b11100100011001101,
    17'b11100010100011111,
    17'b11100001001100110,
    17'b11100000000101001,
    17'b11011111000111101,
    17'b11011101100001010,
    17'b11011100011110110,
    17'b11011011001100110,
    17'b11011011001100110,
    17'b11011100001111011,
    17'b11011100110011010,
    17'b11011101111010111,
    17'b11011111100001010,
    17'b11100111110101110,
    17'b11101001010111000,
    17'b11101010101001000,
    17'b11101100001010010,
    17'b11101101110101110,
    17'b11101110111101100,
    17'b11101111101011100,
    17'b11110000000101001,
    17'b11110000000000000,
    17'b11110000001010010,
    17'b11110000011110110,
    17'b11110000111000011,
    17'b11110001100110011,
    17'b11110010011001101,
    17'b11110100100011111,
    17'b11110110011110110,
    17'b11111000000101001,
    17'b11111001001100110,
    17'b11111001111010111,
    17'b11111001111010111,
    17'b11111001110000101,
    17'b11111010000101001,
    17'b11111001010001111,
    17'b11111000110011010,
    17'b11111000111101100,
    17'b11111001101011100,
    17'b11111001100001010,
    17'b11111001010111000,
    17'b11110100001111011,
    17'b11110010100011111,
    17'b11110001010111000,
    17'b11110000111101100,
    17'b11110000011001101,
    17'b11110000111000011,
    17'b11110000110011010,
    17'b11110001010111000,
    17'b11110000011110110,
    17'b11110000100011111,
    17'b11110000000000000,
    17'b11101111010001111,
    17'b11110001000010100,
    17'b11110011010001111,
    17'b11110100111000011,
    17'b11111001000111101,
    17'b11111010101110001,
    17'b00000100000101001,
    17'b00000101010001111,
    17'b00000111010111000,
    17'b00000110001111011,
    17'b00000011101011100,
    17'b00000110101001000,
    17'b00000101001100110,
    17'b00000100111101100,
    17'b00000110100011111,
    17'b00001000010100100,
    17'b00001000111101100,
    17'b00001011010001111,
    17'b00001100101001000,
    17'b00001100100011111,
    17'b00001010111000011,
    17'b00001001000010100,
    17'b00000111100001010,
    17'b00000110111000011,
    17'b00000011110101110,
    17'b00000010111000011,
    17'b00000111001100110,
    17'b00001000111000011,
    17'b00000111101011100,
    17'b00001001000010100,
    17'b00001101000010100,
    17'b00001100111101100,
    17'b00001110111000011,
    17'b00001111010111000,
    17'b00010001110101110,
    17'b00010011001100110,
    17'b00010011011100001,
    17'b00010101010001111,
    17'b00010100000101001,
    17'b00010010111000011,
    17'b00010001101011100,
    17'b00010011001100110,
    17'b00010110110011010,
    17'b00010110110011010,
    17'b00010101100110011,
    17'b00010100101001000,
    17'b00010100111101100,
    17'b00010010000000000,
    17'b00001011100110011,
    17'b00010100001111011,
    17'b00010101100001010,
    17'b00010110001010010,
    17'b00010100100011111,
    17'b00010111010001111,
    17'b00011000010100100,
    17'b00010010101110001,
    17'b00001110000000000,
    17'b00010000101110001,
    17'b00010000111101100,
    17'b00010000000000000,
    17'b00010001001100110,
    17'b00010100101110001,
    17'b00010100011001101,
    17'b00010101001100110,
    17'b00011101000010100,
    17'b00011100011001101,
    17'b00011010001010010,
    17'b00011010001010010,
    17'b00010101001100110,
    17'b00011010101110001,
    17'b00011000110011010,
    17'b00011101100001010,
    17'b00011101010001111,
    17'b00011100011110110,
    17'b00011100001010010,
    17'b00011010000101001,
    17'b00011101000010100,
    17'b00011010101110001,
    17'b00011001110101110,
    17'b00011001001100110,
    17'b00011010000101001,
    17'b00011010001111011,
    17'b00011001100110011,
    17'b00011001010111000,
    17'b00011001001100110,
    17'b00011000011110110,
    17'b00011000011110110,
    17'b00011001010111000,
    17'b00011001111010111,
    17'b00011001110101110,
    17'b00011001111010111,
    17'b00011001110000101,
    17'b00011001110000101,
    17'b00011001110000101,
    17'b00011001111010111,
    17'b00011001101011100,
    17'b00011001010001111,
    17'b00011000111000011,
    17'b00011000011110110,
    17'b00011001010111000,
    17'b00011010000000000,
    17'b00011010111101100,
    17'b00011011111010111,
    17'b00011100100011111,
    17'b00011100100011111,
    17'b00011100001111011,
    17'b00011100000000000,
    17'b00011011101011100,
    17'b00011011100110011,
    17'b00011011010001111,
    17'b00011011010111000,
    17'b00011011001100110,
    17'b00011010101001000,
    17'b00011010000000000,
    17'b00011001110000101,
    17'b00011001101011100,
    17'b00011000101110001,
    17'b00010111111010111,
    17'b00010110000000000,
    17'b00010101000111101,
    17'b00010011101011100,
    17'b00010101001100110,
    17'b00010110111000011,
    17'b00011001000010100,
    17'b00011000011001101,
    17'b00011000000101001,
    17'b00010111100001010,
    17'b00010111000010100,
    17'b00010110111101100,
    17'b00011000011001101,
    17'b00011000011001101,
    17'b00010110001010010,
    17'b00010101001100110,
    17'b00010100011001101,
    17'b00010011100110011,
    17'b00010010001010010,
    17'b00010001110000101,
    17'b00010000111000011,
    17'b00010000010100100,
    17'b00001111000111101,
    17'b00001110111000011,
    17'b00001110010100100,
    17'b00001101100110011,
    17'b00001101011100001,
    17'b00001101000111101,
    17'b00001100001010010,
    17'b00001011000111101,
    17'b00001010111000011,
    17'b00001011011100001,
    17'b00001011100110011,
    17'b00001011010001111,
    17'b00001011100110011,
    17'b00001011011100001,
    17'b00001010010100100,
    17'b00001010100011111,
    17'b00001011010001111,
    17'b00001100101001000,
    17'b00001110011110110,
    17'b00010000100011111,
    17'b00010001110101110,
    17'b00010001000111101,
    17'b00001111000111101,
    17'b00001101000010100,
    17'b00001010011001101,
    17'b00001000101110001,
    17'b00000111000010100,
    17'b00000101100001010,
    17'b00000100010100100,
    17'b00000100000000000,
    17'b00000100011001101,
    17'b00000100111101100,
    17'b00000110000000000,
    17'b00000110011001101,
    17'b00000110100011111,
    17'b00000110100011111,
    17'b00000110011001101,
    17'b00000110000101001,
    17'b00000101001100110,
    17'b00000100100011111,
    17'b00000100000101001,
    17'b00000011111010111,
    17'b00000011100110011,
    17'b00000011010001111,
    17'b00000011001100110,
    17'b00000011100110011,
    17'b00000100001010010,
    17'b00000100011001101,
    17'b00000100101001000,
    17'b00000100001010010,
    17'b00000011110101110,
    17'b00000011110101110,
    17'b00000011000111101,
    17'b11111101101011100,
    17'b11111110001111011,
    17'b11111110101110001,
    17'b11111111010111000,
    17'b11111111010111000,
    17'b11111111011100001,
    17'b11111111011100001,
    17'b11111110111000011,
    17'b11111110001010010,
    17'b11111101010111000,
    17'b11111100101001000,
    17'b11111011100001010,
    17'b11111010100011111,
    17'b11111001010111000,
    17'b11111000001010010,
    17'b11110111011100001,
    17'b11110111010001111,
    17'b11110111010111000,
    17'b11110111101011100,
    17'b11110111010001111,
    17'b11110110001111011,
    17'b11110100111101100,
    17'b11110010111000011,
    17'b11110001101011100,
    17'b11110000101001000,
    17'b11110000000000000,
    17'b11101110111101100,
    17'b11101110101001000,
    17'b11101110011001101,
    17'b11101110011001101,
    17'b11101110001010010,
    17'b11101110000000000,
    17'b11101110010100100,
    17'b11101110011110110,
    17'b11101111010001111,
    17'b11110000000000000,
    17'b11110000011001101,
    17'b11101111100001010,
    17'b11101110011001101,
    17'b11101101011100001,
    17'b11101100011110110,
    17'b11101011011100001,
    17'b11101010000101001,
    17'b11101000001010010,
    17'b11100101100001010,
    17'b11100011010111000,
    17'b11100010000101001,
    17'b11100010101001000,
    17'b11100010100011111,
    17'b11100001100110011,
    17'b11100000001111011,
    17'b11011111100110011,
    17'b11011110111101100,
    17'b11011111000010100,
    17'b11011110111101100,
    17'b11011110111101100,
    17'b11011111000111101,
    17'b11011111011100001,
    17'b11100000000000000,
    17'b11100000110011010,
    17'b11100010000000000,
    17'b11100001110101110,
    17'b11100001010001111,
    17'b11100000010100100,
    17'b11011111000111101,
    17'b11011110000000000,
    17'b11011100111000011,
    17'b11011100000101001,
    17'b11011011010001111,
    17'b11011010101001000,
    17'b11011001100001010,
    17'b11010111100110011,
    17'b11010101100110011,
    17'b11010100010100100,
    17'b11010100110011010,
    17'b11010100110011010,
    17'b11010011101011100,
    17'b11010010110011010,
    17'b11010010000101001,
    17'b11010010010100100,
    17'b11010011000111101,
    17'b11010010101001000,
    17'b11010001110101110,
    17'b11010001000111101,
    17'b11010001010111000,
    17'b11010001100110011,
    17'b11010001011100001,
    17'b11010000111000011,
    17'b11001111010111000,
    17'b11001101011100001,
    17'b11001100001010010,
    17'b11001011000010100,
    17'b11001011101011100,
    17'b11001101010111000,
    17'b11001100010100100,
    17'b11001010000101001,
    17'b11001001101011100,
    17'b11001110001111011,
    17'b11001110011110110,
    17'b11001110000101001,
    17'b11001110001111011,
    17'b11001110000000000,
    17'b11001101000010100,
    17'b11001110000101001,
    17'b11001111100110011,
    17'b11001111001100110,
    17'b11001110100011111,
    17'b11001101010111000,
    17'b11001100000101001,
    17'b11001010101110001,
    17'b11001010001111011,
    17'b11001001110101110,
    17'b11001001101011100,
    17'b11001010001010010,
    17'b11001010101110001,
    17'b11001011010001111,
    17'b11001010010100100,
    17'b11001011010001111,
    17'b11001110101001000,
    17'b11010000111101100,
    17'b11010001010111000,
    17'b11010000011001101,
    17'b11001101011100001,
    17'b11001100000101001,
    17'b11001100111000011,
    17'b11001110100011111,
    17'b11010001010111000,
    17'b11010010101001000,
    17'b11010011001100110,
    17'b11010011100110011,
    17'b11010011111010111,
    17'b11010100011110110,
    17'b11010100011110110,
    17'b11010100000101001,
    17'b11010011110000101,
    17'b11010011111010111,
    17'b11010011100110011,
    17'b11010011000111101,
    17'b11010010100011111,
    17'b11010001100001010,
    17'b11010000001010010,
    17'b11001111000111101,
    17'b11001110011001101,
    17'b11001101100110011,
    17'b11001110111000011,
    17'b11001111010001111,
    17'b11010000001010010,
    17'b11010000111101100,
    17'b11010010111000011,
    17'b11010011110101110,
    17'b11010101010001111,
    17'b11010110101001000,
    17'b11011001000010100,
    17'b11011110011001101,
    17'b11100000101110001,
    17'b11100001110101110,
    17'b11100001111010111,
    17'b11100000110011010,
    17'b11100001011100001,
    17'b11100001011100001,
    17'b11100010001010010,
    17'b11100011001100110,
    17'b11100010000101001,
    17'b11100010011110110,
    17'b11100010110011010,
    17'b11100001010111000,
    17'b11011111000111101,
    17'b11011110111101100,
    17'b11011111001100110,
    17'b11011110011001101,
    17'b11011101011100001,
    17'b11011101111010111,
    17'b11011101110101110,
    17'b11011101111010111,
    17'b11011110001010010,
    17'b11011110011001101,
    17'b11011111111010111,
    17'b11100000111000011,
    17'b11100010011001101,
    17'b11100011001100110,
    17'b11100011100110011,
    17'b11100100010100100,
    17'b11100100110011010,
    17'b11100110110011010,
    17'b11101000010100100,
    17'b11101010010100100,
    17'b11101010101001000,
    17'b11101010001111011,
    17'b11101100011001101,
    17'b11101110100011111,
    17'b11110000011001101,
    17'b11110001101011100,
    17'b11110001011100001,
    17'b11110001010001111,
    17'b11110000111101100,
    17'b11110000111101100,
    17'b11110001001100110,
    17'b11110000111000011,
    17'b11110000011110110,
    17'b11101111100110011,
    17'b11101111001100110,
    17'b11101110111101100,
    17'b11101111110000101,
    17'b11110000011001101,
    17'b11110000110011010,
    17'b11110010111101100,
    17'b11110011010111000,
    17'b11110011011100001,
    17'b11110011010001111,
    17'b11110100110011010,
    17'b11110110010100100,
    17'b11110110101110001,
    17'b11110111000111101,
    17'b11110110101001000,
    17'b11110110011001101,
    17'b11110110111000011,
    17'b11110111100110011,
    17'b11111001001100110,
    17'b11111010001111011,
    17'b11111011101011100,
    17'b11111100110011010,
    17'b11111110001111011,
    17'b11111111000111101,
    17'b00000000001010010,
    17'b00000000100011111,
    17'b00000000011001101,
    17'b00000000011110110,
    17'b00000001000111101,
    17'b00000010010100100,
    17'b00000011100110011,
    17'b00000101010001111,
    17'b00000111010001111,
    17'b00000111110000101,
    17'b00001000111101100,
    17'b00001010001010010,
    17'b00001010010100100,
    17'b00001010100011111,
    17'b00001010011001101,
    17'b00001011001100110,
    17'b00001011111010111,
    17'b00001101000010100,
    17'b00001110111101100,
    17'b00001011001100110,
    17'b00001010000000000,
    17'b00001001101011100,
    17'b00000110101001000,
    17'b00000101111010111,
    17'b00001000101110001,
    17'b00001011101011100,
    17'b00001101010111000,
    17'b00001110101110001,
    17'b00001111001100110,
    17'b00001111010001111,
    17'b00001111111010111,
    17'b00001100110011010,
    17'b00001100011110110,
    17'b00001011100001010,
    17'b00001010111101100,
    17'b00001100101001000,
    17'b00001101101011100,
    17'b00001110101001000,
    17'b00010000000000000,
    17'b00010001111010111,
    17'b00010011001100110,
    17'b00010011111010111,
    17'b00010100010100100,
    17'b00010100111000011,
    17'b00010101111010111,
    17'b00010110110011010,
    17'b00010111110000101,
    17'b00011000010100100,
    17'b00011000110011010,
    17'b00011001011100001,
    17'b00011001100001010,
    17'b00011010001111011,
    17'b00011010110011010,
    17'b00011010101110001,
    17'b00011010011001101,
    17'b00011010011001101,
    17'b00011010011001101,
    17'b00011011000111101,
    17'b00011100000101001,
    17'b00011100111000011,
    17'b00011111011100001,
    17'b00100011101011100,
    17'b00100111000111101,
    17'b00100110111000011,
    17'b00100101001100110,
    17'b00100011000010100,
    17'b00100000111101100,
    17'b00011100110011010,
    17'b00011100011001101,
    17'b00011100000101001,
    17'b00011100010100100,
    17'b00011100010100100,
    17'b00011101010001111,
    17'b00011101111010111,
    17'b00011101110000101,
    17'b00011110001111011,
    17'b00011111000111101,
    17'b00011110110011010,
    17'b00011110001010010,
    17'b00011101101011100,
    17'b00011100111000011,
    17'b00011100111000011,
    17'b00011011110101110,
    17'b00011011010001111,
    17'b00011011101011100,
    17'b00011100001010010,
    17'b00011101001100110,
    17'b00011110001111011,
    17'b00011111001100110,
    17'b00011111001100110,
    17'b00011111110101110,
    17'b00100000000000000,
    17'b00100000000000000,
    17'b00100000101110001,
    17'b00100001100110011,
    17'b00100001110000101,
    17'b00100010001111011,
    17'b00100011010001111,
    17'b00100011101011100,
    17'b00100100010100100,
    17'b00100101100001010,
    17'b00100101110101110,
    17'b00100100100011111,
    17'b00100010100011111,
    17'b00100000110011010,
    17'b00011111001100110,
    17'b00011011000111101,
    17'b00011011001100110,
    17'b00011010101001000,
    17'b00011010011110110,
    17'b00011001110000101,
    17'b00011000100011111,
    17'b00010110011110110,
    17'b00010011010111000,
    17'b00010001111010111,
    17'b00010000111000011,
    17'b00010000011001101,
    17'b00001110101001000,
    17'b00001101111010111,
    17'b00001101101011100,
    17'b00001110000000000,
    17'b00001110000000000,
    17'b00001110000000000,
    17'b00001110001111011,
    17'b00001101010111000,
    17'b00001101000010100,
    17'b00001100111000011,
    17'b00001100000000000,
    17'b00001010011110110,
    17'b00001010000000000,
    17'b00001001011100001,
    17'b00000111111010111,
    17'b00000111100001010,
    17'b00000111010001111,
    17'b00000111010001111,
    17'b00000100111000011,
    17'b00000000001010010,
    17'b11111101111010111,
    17'b11111011110000101,
    17'b11111001111010111,
    17'b11111010111000011,
    17'b11111100011110110,
    17'b11111100000101001,
    17'b11111000010100100,
    17'b11110011000111101,
    17'b11110001100110011,
    17'b11110100101001000,
    17'b11110111000010100,
    17'b11110111000010100,
    17'b11110111000111101,
    17'b11110111000010100,
    17'b11110110000101001,
    17'b11110011001100110,
    17'b11110011000010100,
    17'b11110101100110011,
    17'b11110110100011111,
    17'b11110110111101100,
    17'b11110111100110011,
    17'b11110111010111000,
    17'b11110110011001101,
    17'b11110100101001000,
    17'b11101110010100100,
    17'b11101100110011010,
    17'b11101011110101110,
    17'b11101001101011100,
    17'b11100111111010111,
    17'b11100100100011111,
    17'b11100010011001101,
    17'b11100111000111101,
    17'b11101000011001101,
    17'b11101000010100100,
    17'b11100111100001010,
    17'b11100101011100001,
    17'b11100001000010100,
    17'b11100100111000011,
    17'b11100101010001111,
    17'b11100100000000000,
    17'b11100011010001111,
    17'b11100011001100110,
    17'b11011110001111011,
    17'b11100010001010010,
    17'b11100101110000101,
    17'b11100101011100001,
    17'b11100101010111000,
    17'b11100110001111011,
    17'b11100110101110001,
    17'b11100101110000101,
    17'b11100101000010100,
    17'b11100100011110110,
    17'b11100011110101110,
    17'b11100011000111101,
    17'b11100101110000101,
    17'b11100110100011111,
    17'b11100111000010100,
    17'b11100110000000000,
    17'b11100100111000011,
    17'b11100010110011010,
    17'b11100001100001010,
    17'b11100000010100100,
    17'b11011111110101110,
    17'b11011111110101110,
    17'b11100000011001101,
    17'b11100001100001010,
    17'b11100010001010010,
    17'b11100010000101001,
    17'b11100001010001111,
    17'b11100000111101100,
    17'b11100000100011111,
    17'b11100000001010010,
    17'b11011111100110011,
    17'b11011111100001010,
    17'b11100000000000000,
    17'b11100001001100110,
    17'b11100001100110011,
    17'b11100001010001111,
    17'b11100001001100110,
    17'b11100001000010100,
    17'b11100000101001000,
    17'b11011110111000011,
    17'b11011100101001000,
    17'b11011011010111000,
    17'b11011010101001000,
    17'b11011010101001000,
    17'b11011010000101001,
    17'b11011001001100110,
    17'b11010111110101110,
    17'b11010001011100001,
    17'b11010000110011010,
    17'b11010000000101001,
    17'b11010000011001101,
    17'b11010000100011111,
    17'b11010000011001101,
    17'b11010000101001000,
    17'b11010001110101110,
    17'b11010011001100110,
    17'b11010100010100100,
    17'b11010100101110001,
    17'b11010100110011010,
    17'b11010100110011010,
    17'b11010101000111101,
    17'b11010101100001010,
    17'b11010110001010010,
    17'b11010110001111011,
    17'b11010110011110110,
    17'b11010110101110001,
    17'b11010111010001111,
    17'b11010111000111101,
    17'b11010110101110001,
    17'b11010101100001010,
    17'b11010100101001000,
    17'b11010011100110011,
    17'b11010010101001000,
    17'b11010001101011100,
    17'b11010001000111101,
    17'b11010000110011010,
    17'b11010000000101001,
    17'b11001111001100110,
    17'b11001110010100100,
    17'b11001101010001111,
    17'b11001100011110110,
    17'b11001011010111000,
    17'b11001010111101100,
    17'b11001010001111011,
    17'b11001010000101001,
    17'b11001000101110001,
    17'b11000111111010111,
    17'b11001000001010010,
    17'b11001000110011010,
    17'b11001111010001111,
    17'b11001111100001010,
    17'b11001111000111101,
    17'b11001110011001101,
    17'b11001110011001101,
    17'b11001110001111011,
    17'b11001110001010010,
    17'b11001101110101110,
    17'b11001100110011010,
    17'b11001101010001111,
    17'b11001100000101001,
    17'b11001011000010100,
    17'b11001010111000011,
    17'b11001001100001010,
    17'b11001000110011010,
    17'b11000111100110011,
    17'b11000110101001000,
    17'b11000101011100001,
    17'b11000100100011111,
    17'b11000100000101001,
    17'b11000010000101001,
    17'b11000000110011010,
    17'b10111111100001010,
    17'b11000000011110110,
    17'b11000000111000011,
    17'b10111111101011100,
    17'b11000011000010100,
    17'b11000011100001010,
    17'b11000101000111101,
    17'b11001101110000101,
    17'b11010100101001000,
    17'b11001100011110110,
    17'b11000110101110001,
    17'b10111100011001101,
    17'b10110111110101110,
    17'b10110101110101110,
    17'b10110101100001010,
    17'b10111100001111011,
    17'b10111101000111101,
    17'b11000001010111000,
    17'b11000001000010100,
    17'b11000000111000011,
    17'b10111110100011111,
    17'b10111100000101001,
    17'b10111010000101001,
    17'b10111001100001010,
    17'b10111010001010010,
    17'b10111010010100100,
    17'b10111010001111011,
    17'b10111001110101110,
    17'b10111001110101110,
    17'b10111010001010010,
    17'b10111010111101100,
    17'b10111011010111000,
    17'b10111100000000000,
    17'b10111011101011100,
    17'b10111101010111000,
    17'b10111110000000000,
    17'b10111111010111000,
    17'b10111111010001111,
    17'b11000001111010111,
    17'b11000001111010111,
    17'b11000010000000000,
    17'b11000000001111011,
    17'b11000000001111011,
    17'b10111110001010010,
    17'b10111100001111011,
    17'b10111110001111011,
    17'b10111100011001101,
    17'b10111000011110110,
    17'b10111100101001000,
    17'b10111100001111011,
    17'b10110001000111101,
    17'b11000010110011010,
    17'b11000101001100110,
    17'b11000101110101110,
    17'b11000100011001101,
    17'b11000100000101001,
    17'b11000010111000011,
    17'b11000000001010010,
    17'b10111101011100001,
    17'b10111011110101110,
    17'b10111100011001101,
    17'b10111101000010100,
    17'b10111101001100110,
    17'b10111101110101110,
    17'b10111110011001101,
    17'b10111110111101100,
    17'b10111111101011100,
    17'b11000000001010010,
    17'b11000000100011111,
    17'b11000001000111101,
    17'b11000001100001010,
    17'b11000001110101110,
    17'b11000010000101001,
    17'b11000010111101100,
    17'b11000011000111101,
    17'b11000010011110110,
    17'b11000011000010100,
    17'b11000100101110001,
    17'b11000010000000000,
    17'b11000100011001101,
    17'b11000010000101001,
    17'b10111110010100100,
    17'b10111101010111000,
    17'b10111101101011100,
    17'b10111110111101100,
    17'b10111111011100001,
    17'b10111110101001000,
    17'b10111110000000000,
    17'b10111110010100100,
    17'b10111110001111011,
    17'b10111101110101110,
    17'b10111110001010010,
    17'b10111111010111000,
    17'b10111110100011111,
    17'b10111111010001111,
    17'b10111111110000101,
    17'b11000001000111101,
    17'b11000001000010100,
    17'b10111111111010111,
    17'b10111111110101110,
    17'b11000001011100001,
    17'b11000000110011010,
    17'b10111110101001000,
    17'b10111101101011100,
    17'b10111110001111011,
    17'b10111011010111000,
    17'b10111100110011010,
    17'b10111100000101001,
    17'b10111010111101100,
    17'b10111100001111011,
    17'b10111111001100110,
    17'b10111111100001010,
    17'b10111111010111000,
    17'b11000000010100100,
    17'b11000011000111101,
    17'b11000110001111011,
    17'b11001011110000101,
    17'b11001010011001101,
    17'b11001110011110110,
    17'b11001111111010111,
    17'b11001111000010100,
    17'b11010001000111101,
    17'b11010000111101100,
    17'b11010001000010100,
    17'b11010000101110001,
    17'b11010000111000011,
    17'b11010000111101100,
    17'b11010000011001101,
    17'b11001111101011100,
    17'b11001111010001111,
    17'b11001110010100100,
    17'b11001111001100110,
    17'b11010000100011111,
    17'b11010001110101110,
    17'b11010100000000000,
    17'b11010101000010100,
    17'b11010101111010111,
    17'b11010110111101100,
    17'b11011000011001101,
    17'b11011000101110001,
    17'b11011000111101100,
    17'b11011001011100001,
    17'b11011001100110011,
    17'b11011010000101001,
    17'b11011010111101100,
    17'b11011100000101001,
    17'b11011100110011010,
    17'b11011101011100001,
    17'b11011101100110011,
    17'b11011101100001010,
    17'b11011101100110011,
    17'b11011101101011100,
    17'b11011101110000101,
    17'b11011010101110001,
    17'b11011011000010100,
    17'b11011011100001010,
    17'b11011011111010111,
    17'b11011100011001101,
    17'b11011101000111101,
    17'b11011101110101110,
    17'b11011110111101100,
    17'b11100000000101001,
    17'b11100000110011010,
    17'b11011111110000101,
    17'b11011111000010100,
    17'b11011110011110110,
    17'b11011110001010010,
    17'b11011110011110110,
    17'b11011111000010100,
    17'b11100000001010010,
    17'b11100010000101001,
    17'b11100100000101001,
    17'b11100101111010111,
    17'b11100111110000101,
    17'b11101001000010100,
    17'b11101010100011111,
    17'b11101011010001111,
    17'b11101001110101110,
    17'b11101010000000000,
    17'b11101010110011010,
    17'b11101010111101100,
    17'b11101000111101100,
    17'b11101000110011010,
    17'b11101000110011010,
    17'b11100101011100001,
    17'b11100100001111011,
    17'b11100010111000011,
    17'b11100001001100110,
    17'b11011111011100001,
    17'b11011110100011111,
    17'b11011110000101001,
    17'b11011101001100110,
    17'b11011100000101001,
    17'b11011101110101110,
    17'b11011110111101100,
    17'b11011111010111000,
    17'b11011111001100110,
    17'b11011111100110011,
    17'b11100000111101100,
    17'b11100011110000101,
    17'b11100101010111000,
    17'b11100110101001000,
    17'b11100110111000011,
    17'b11101000101001000,
    17'b11101010011001101,
    17'b11101010001010010,
    17'b11101010111000011,
    17'b11101110011110110,
    17'b11110001011100001,
    17'b11110010111000011,
    17'b11110010101001000,
    17'b11110010010100100,
    17'b11110001110000101,
    17'b11110000110011010,
    17'b11110000011110110,
    17'b11101111101011100,
    17'b11110000001010010,
    17'b11110001010001111,
    17'b11110001110000101,
    17'b11110001100110011,
    17'b11110001111010111,
    17'b11110001101011100,
    17'b11110010000000000,
    17'b11110001111010111,
    17'b11110010000101001,
    17'b11110001110101110,
    17'b11110001010001111,
    17'b11110000100011111,
    17'b11110000010100100,
    17'b11110000101110001,
    17'b11110000000101001,
    17'b11101111111010111,
    17'b11110001001100110,
    17'b11110010111000011,
    17'b11110100001010010,
    17'b11110100011110110,
    17'b11110101000111101,
    17'b11110110001010010,
    17'b11111000010100100,
    17'b11111011101011100,
    17'b11111100000101001,
    17'b11111100000101001,
    17'b11111100001010010,
    17'b11111011100001010,
    17'b11111010101001000,
    17'b11111001100001010,
    17'b11111000111101100,
    17'b11111000100011111,
    17'b11111000000000000,
    17'b11110111111010111,
    17'b11111000000101001,
    17'b11111000110011010,
    17'b11111001011100001,
    17'b11111001011100001,
    17'b11111001000010100,
    17'b11111000111000011,
    17'b11111000111000011,
    17'b11111000111000011,
    17'b11111000101110001,
    17'b11111000101110001,
    17'b11111001010111000,
    17'b11111001101011100,
    17'b11111001111010111,
    17'b11111000111000011,
    17'b11111100010100100,
    17'b11111101000111101,
    17'b11111101101011100,
    17'b11111101000111101,
    17'b11111100011001101,
    17'b11111011101011100,
    17'b11111011010111000,
    17'b11111011010001111,
    17'b11111011010001111,
    17'b11111011011100001,
    17'b11111010101110001,
    17'b11111010011110110,
    17'b11111010000101001,
    17'b11111010000000000,
    17'b11111001011100001,
    17'b11111000111101100,
    17'b11110111111010111,
    17'b11111010000101001,
    17'b11111010111000011,
    17'b11111000000000000,
    17'b11111010001111011,
    17'b11111001101011100,
    17'b11111000000101001,
    17'b11110101010001111,
    17'b11110000101001000,
    17'b11101101100001010,
    17'b11101011000111101,
    17'b11101001110101110,
    17'b11101000101001000,
    17'b11101000100011111,
    17'b11100111100001010,
    17'b11100110000000000,
    17'b11100001100001010,
    17'b11011110100011111,
    17'b11011011110000101,
    17'b11011010101110001,
    17'b11011010101110001,
    17'b11011100011001101,
    17'b11011010001010010,
    17'b11011001010001111,
    17'b11011010110011010,
    17'b11011010011110110,
    17'b11011001100001010,
    17'b11010111110000101,
    17'b11010101100001010,
    17'b11010011110000101,
    17'b11010011010001111,
    17'b11010011000111101,
    17'b11010011100110011,
    17'b11010011010111000,
    17'b11010011011100001,
    17'b11010011000010100,
    17'b11010010111101100,
    17'b11010010011110110,
    17'b11010010000101001,
    17'b11010010010100100,
    17'b11010000111000011,
    17'b11001101010111000,
    17'b11001010000000000,
    17'b11001001100110011,
    17'b11001010000000000,
    17'b11001011001100110,
    17'b11010000000000000,
    17'b11011001100001010,
    17'b11010111011100001,
    17'b11010101110101110,
    17'b11010010111000011,
    17'b11001100100011111,
    17'b11001000001010010,
    17'b11000100111101100,
    17'b11000011110000101,
    17'b11000011010111000,
    17'b11000011101011100,
    17'b11000011011100001,
    17'b11000011100001010,
    17'b11000011110000101,
    17'b11000100101110001,
    17'b11000110000000000,
    17'b11001000100011111,
    17'b11001010101110001,
    17'b11001100101110001,
    17'b11001111000111101,
    17'b11010000101001000,
    17'b11010010000000000,
    17'b11010010111000011,
    17'b11010100000000000,
    17'b11010011100001010,
    17'b11010011001100110,
    17'b11010010011001101,
    17'b11010010000101001,
    17'b11010001100110011,
    17'b11010001100001010,
    17'b11010001010001111,
    17'b11010000111101100,
    17'b11001111110101110,
    17'b11001000001111011,
    17'b11001000101001000,
    17'b11001001000010100,
    17'b11001011100001010,
    17'b11001110101001000,
    17'b11010010011110110,
    17'b11010100010100100,
    17'b11010101111010111,
    17'b11010110001010010,
    17'b11010101100001010,
    17'b11010011110101110,
    17'b11010011001100110,
    17'b11010010101110001,
    17'b11010010011110110,
    17'b11010011000111101,
    17'b11010100011001101,
    17'b11010110100011111,
    17'b11011000001111011,
    17'b11011001101011100,
    17'b11011001100001010,
    17'b11011010100011111,
    17'b11011001110101110,
    17'b11011010000101001,
    17'b11011000011001101,
    17'b11010111010111000,
    17'b11011001001100110,
    17'b11011110101110001,
    17'b11100011011100001,
    17'b11011111110101110,
    17'b11100001110000101,
    17'b11100010111101100,
    17'b11100101011100001,
    17'b11100101010001111,
    17'b11100011000111101,
    17'b11011110110011010,
    17'b11011010011110110,
    17'b11010101111010111,
    17'b11010100001010010,
    17'b11010010101110001,
    17'b11010011000010100,
    17'b11010011100001010,
    17'b11010011110000101,
    17'b11010100011001101,
    17'b11010101010001111,
    17'b11010110100011111,
    17'b11010111110101110,
    17'b11011001111010111,
    17'b11011010110011010,
    17'b11011011000111101,
    17'b11011011010111000,
    17'b11011011111010111,
    17'b11011101011100001,
    17'b11100000111000011,
    17'b11100010001111011,
    17'b11100011010001111,
    17'b11100100011001101,
    17'b11100101110000101,
    17'b11100111110101110,
    17'b11101000011110110,
    17'b11101001100110011,
    17'b11101010011110110,
    17'b11101010111000011,
    17'b11101010000000000,
    17'b11101000001010010,
    17'b11100101000010100,
    17'b11100010000000000,
    17'b11011111010001111,
    17'b11011100101110001,
    17'b11011001110101110,
    17'b11010111110101110,
    17'b11010110010100100,
    17'b11010101000010100,
    17'b11010100101001000,
    17'b11010101011100001,
    17'b11010110001010010,
    17'b11010110110011010,
    17'b11010111000111101,
    17'b11010111110101110,
    17'b11011000010100100,
    17'b11011000000101001,
    17'b11010111101011100,
    17'b11010111011100001,
    17'b11010111010111000,
    17'b11010111000111101,
    17'b11010110110011010,
    17'b11010110110011010,
    17'b11010110111000011,
    17'b11010110001111011,
    17'b11010110001010010,
    17'b11010101100001010,
    17'b11010010110011010,
    17'b11010010011001101,
    17'b11010000010100100,
    17'b11001110000000000,
    17'b11001100100011111,
    17'b11001100001111011,
    17'b11001100011001101,
    17'b11001100000000000,
    17'b11001010110011010,
    17'b11001001000111101,
    17'b11000111100110011,
    17'b11000111100110011,
    17'b11001000010100100,
    17'b11001001011100001,
    17'b11001010101110001,
    17'b11001011011100001,
    17'b11001011000111101,
    17'b11001010011110110,
    17'b11001001010001111,
    17'b11001000001010010,
    17'b11000111010001111,
    17'b11000110111000011,
    17'b11000110110011010,
    17'b11000110001111011,
    17'b11000110000101001,
    17'b11001001111010111,
    17'b11001001101011100,
    17'b11000111010111000,
    17'b11000101000010100,
    17'b11000010001010010,
    17'b10111111111010111,
    17'b10111110001010010,
    17'b10111101110101110,
    17'b10111110011110110,
    17'b10111110111101100,
    17'b10111111110000101,
    17'b11000000000101001,
    17'b11000000110011010,
    17'b11000001000111101,
    17'b11000000111101100,
    17'b11000000011001101,
    17'b10111111100001010,
    17'b10111110100011111,
    17'b10111110010100100,
    17'b10111110000000000,
    17'b10111101100110011,
    17'b10111101000010100,
    17'b10111100100011111,
    17'b10111011101011100,
    17'b10111011010001111,
    17'b10111010101110001,
    17'b10111000110011010,
    17'b10110110111101100,
    17'b10110100001010010,
    17'b10110101100001010,
    17'b10110110110011010,
    17'b10110110100011111,
    17'b10110110111000011,
    17'b10111001001100110,
    17'b10111011000010100,
    17'b10111100111000011,
    17'b10111110110011010,
    17'b11000000101110001,
    17'b11000001100110011,
    17'b11000001110101110,
    17'b11000010000000000,
    17'b11000001011100001,
    17'b11000001001100110,
    17'b11000001100110011,
    17'b11000010011001101,
    17'b11000011110000101,
    17'b11000100011110110,
    17'b11000101001100110,
    17'b11000101100001010,
    17'b11000110001010010,
    17'b11000110101001000,
    17'b11000111001100110,
    17'b11000111010001111,
    17'b11000111010111000,
    17'b11000111101011100,
    17'b11000111111010111,
    17'b11001000011110110,
    17'b11001000110011010,
    17'b11001010000000000,
    17'b11001010110011010,
    17'b11001011100110011,
    17'b11001100000101001,
    17'b11001100011110110,
    17'b11001101000010100,
    17'b11001101101011100,
    17'b11001110111000011,
    17'b11010000001111011,
    17'b11010001110101110,
    17'b11010011000010100,
    17'b11010100101001000,
    17'b11010101110000101,
    17'b11010111011100001,
    17'b11011000111101100,
    17'b11011010001010010,
    17'b11011010111000011,
    17'b11011011010111000,
    17'b11011100000101001,
    17'b11011100010100100,
    17'b11011101001100110,
    17'b11011110010100100,
    17'b11011111110000101,
    17'b11100000001111011,
    17'b11100000011001101
};

parameter logic signed [`ACC_WIDTH-1:0] AY_TEST_VECTOR[`NUM_ELEMENTS] = {
    17'b00101001010001111,
    17'b00101001000111101,
    17'b00101000101110001,
    17'b00101000001010010,
    17'b00100111101011100,
    17'b00100110101110001,
    17'b00100110001111011,
    17'b00100101110000101,
    17'b00100101001100110,
    17'b00100011111010111,
    17'b00100010101001000,
    17'b00100001110000101,
    17'b00100001011100001,
    17'b00100001011100001,
    17'b00100001010001111,
    17'b00100001000111101,
    17'b00100000100011111,
    17'b00011111110101110,
    17'b00011111010001111,
    17'b00011110100011111,
    17'b00011110000000000,
    17'b00011100111101100,
    17'b00011100001111011,
    17'b00011011100110011,
    17'b00011011000111101,
    17'b00011010010100100,
    17'b00011001101011100,
    17'b00011000111101100,
    17'b00011000001010010,
    17'b00010110101001000,
    17'b00010101001100110,
    17'b00010011110000101,
    17'b00010001110000101,
    17'b00010000000101001,
    17'b00001110111000011,
    17'b00001101010001111,
    17'b00001010101110001,
    17'b00001001110101110,
    17'b00001001101011100,
    17'b00001010001010010,
    17'b00001010011001101,
    17'b00001001101011100,
    17'b00001000010100100,
    17'b00000110111000011,
    17'b00000101110101110,
    17'b00000101010001111,
    17'b00000100111101100,
    17'b00000100011110110,
    17'b00000011100001010,
    17'b00000010011001101,
    17'b00000001010111000,
    17'b00000000101110001,
    17'b11111111110101110,
    17'b11111111010001111,
    17'b11111110101110001,
    17'b11111110000101001,
    17'b11111101110000101,
    17'b11111101100110011,
    17'b11111101100001010,
    17'b11111101100110011,
    17'b11111101110101110,
    17'b11111110000000000,
    17'b11111110001111011,
    17'b11111110001111011,
    17'b11111100011001101,
    17'b11111010011110110,
    17'b11111010001010010,
    17'b11111010111101100,
    17'b11111011100001010,
    17'b11111100011110110,
    17'b11111110000000000,
    17'b11111111101011100,
    17'b00000001010111000,
    17'b00000010011110110,
    17'b00000100000000000,
    17'b00001001101011100,
    17'b00010010000000000,
    17'b00010110001010010,
    17'b00011011100110011,
    17'b00100001100110011,
    17'b00100110101001000,
    17'b00011110001111011,
    17'b00001100101110001,
    17'b11111001101011100,
    17'b11101100101001000,
    17'b11101011000010100,
    17'b11110100011001101,
    17'b11111110001010010,
    17'b00000010110011010,
    17'b00000011000111101,
    17'b00000010111000011,
    17'b00000100000101001,
    17'b00000110000101001,
    17'b00000111010001111,
    17'b00000101010001111,
    17'b00000001110000101,
    17'b11111101111010111,
    17'b11111011010001111,
    17'b11111100000000000,
    17'b11111101000111101,
    17'b11111101010111000,
    17'b11111110110011010,
    17'b00000000111000011,
    17'b00000100011001101,
    17'b00000111100001010,
    17'b00001010010100100,
    17'b00001111000010100,
    17'b00010001000010100,
    17'b00010001110101110,
    17'b00010011000111101,
    17'b00010011000010100,
    17'b00010000000101001,
    17'b00001101000010100,
    17'b00001011010111000,
    17'b00001011010111000,
    17'b00001100010100100,
    17'b00001100111000011,
    17'b00001101000111101,
    17'b00001101010111000,
    17'b00001101100110011,
    17'b00001101110000101,
    17'b00010001111010111,
    17'b00010110001111011,
    17'b00010000110011010,
    17'b00001011101011100,
    17'b00001011110000101,
    17'b00001010110011010,
    17'b00001010110011010,
    17'b00001100111101100,
    17'b00001101110000101,
    17'b00001110000000000,
    17'b00001101111010111,
    17'b00001100011001101,
    17'b00001100010100100,
    17'b00001100000000000,
    17'b00001011000111101,
    17'b00001100000101001,
    17'b00001101110000101,
    17'b00001100011110110,
    17'b00001011110000101,
    17'b00000111110000101,
    17'b00000100010100100,
    17'b00000001010111000,
    17'b00000001010111000,
    17'b00000001100110011,
    17'b00000010011001101,
    17'b00000010111101100,
    17'b00000011110000101,
    17'b00001000001010010,
    17'b00001001100001010,
    17'b00001010000000000,
    17'b00001010000101001,
    17'b00000111110000101,
    17'b00000110011001101,
    17'b00000101100001010,
    17'b00000101000010100,
    17'b00000111100110011,
    17'b00001011011100001,
    17'b00001111011100001,
    17'b00010010001010010,
    17'b00010010101110001,
    17'b00010001011100001,
    17'b00010000000101001,
    17'b00001111001100110,
    17'b00001101010111000,
    17'b00001100011110110,
    17'b00001011010001111,
    17'b00001100101001000,
    17'b00001101100110011,
    17'b00001010101110001,
    17'b00000111000010100,
    17'b00000100001111011,
    17'b00000010001111011,
    17'b00000000110011010,
    17'b11111110111101100,
    17'b11111101000111101,
    17'b11111010111000011,
    17'b11111010110011010,
    17'b11111100100011111,
    17'b11111010000101001,
    17'b11110101110000101,
    17'b11110100110011010,
    17'b11111001100001010,
    17'b00000010101001000,
    17'b00001010100011111,
    17'b00010010111000011,
    17'b00011010100011111,
    17'b00100000100011111,
    17'b00100100101110001,
    17'b00100100001111011,
    17'b00100011000010100,
    17'b00100010011110110,
    17'b00100001000111101,
    17'b00011110011001101,
    17'b00011001000111101,
    17'b00010001111010111,
    17'b00000110001111011,
    17'b11111101100110011,
    17'b11110101010111000,
    17'b11101110011110110,
    17'b11100110000101001,
    17'b11011110101110001,
    17'b11011100101110001,
    17'b11011100101001000,
    17'b11011001110101110,
    17'b11010111100110011,
    17'b11011000111101100,
    17'b11011001100001010,
    17'b11011100101001000,
    17'b11100000111000011,
    17'b11100101010001111,
    17'b11101001010001111,
    17'b11101100111000011,
    17'b11110000001111011,
    17'b11110001110101110,
    17'b11110010111101100,
    17'b11110100000000000,
    17'b11110110011001101,
    17'b11111001000010100,
    17'b11111100001111011,
    17'b11111111101011100,
    17'b00000011110000101,
    17'b00000101110000101,
    17'b00000110001111011,
    17'b00000101001100110,
    17'b00000010111000011,
    17'b11111111000010100,
    17'b11111100001111011,
    17'b11111010001010010,
    17'b11111000110011010,
    17'b11111000010100100,
    17'b11111000101110001,
    17'b11111001011100001,
    17'b11111010010100100,
    17'b11111011010001111,
    17'b11111100000101001,
    17'b11111100110011010,
    17'b11111101100110011,
    17'b11111110001111011,
    17'b11111110111101100,
    17'b11111111110101110,
    17'b00000010001010010,
    17'b00000100100011111,
    17'b00000111010111000,
    17'b00001010000000000,
    17'b00001010111000011,
    17'b00001000111000011,
    17'b00000101111010111,
    17'b11111100110011010,
    17'b00000101101011100,
    17'b00000111010111000,
    17'b00001011100001010,
    17'b00001001010111000,
    17'b00001010111101100,
    17'b00001000100011111,
    17'b00001011010001111,
    17'b00001101100001010,
    17'b00001011010001111,
    17'b00000010001111011,
    17'b11111010101001000,
    17'b11110000011110110,
    17'b11101000110011010,
    17'b11100010111000011,
    17'b11100011101011100,
    17'b11100111001100110,
    17'b11101010001010010,
    17'b11101011010111000,
    17'b11101010101001000,
    17'b11101000111000011,
    17'b11100111000010100,
    17'b11100101110000101,
    17'b11100010110011010,
    17'b11100001010111000,
    17'b11100001000010100,
    17'b11100001110101110,
    17'b11100010110011010,
    17'b11100100010100100,
    17'b11100110001111011,
    17'b11100111000010100,
    17'b11100111110101110,
    17'b11101000010100100,
    17'b11101001000111101,
    17'b11101001111010111,
    17'b11101100100011111,
    17'b11110001100001010,
    17'b11110101010001111,
    17'b11110111101011100,
    17'b11111010011110110,
    17'b11111011101011100,
    17'b11111100011001101,
    17'b11111100110011010,
    17'b11111101000010100,
    17'b11111101000010100,
    17'b11111101010111000,
    17'b11111101010111000,
    17'b11111101001100110,
    17'b11111101010001111,
    17'b11111101001100110,
    17'b11111101010001111,
    17'b11111101000111101,
    17'b11111101010001111,
    17'b11111101001100110,
    17'b11111101010001111,
    17'b11111101010001111,
    17'b11111101010001111,
    17'b11111101010111000,
    17'b11111101011100001,
    17'b11111101100001010,
    17'b11111101100001010,
    17'b11111101100110011,
    17'b11111101100001010,
    17'b11111101011100001,
    17'b11111101100001010,
    17'b11111101100001010,
    17'b11111101100110011,
    17'b11111101100110011,
    17'b11111101100001010,
    17'b11111101100001010,
    17'b11111101100110011,
    17'b11111101011100001,
    17'b11111101010111000,
    17'b11111101010111000,
    17'b11111101010111000,
    17'b11111101010111000,
    17'b11111101010001111,
    17'b11111101010111000,
    17'b11111101010001111,
    17'b11111101010001111,
    17'b11111101010111000,
    17'b11111101010111000,
    17'b11111101010111000,
    17'b11111101011100001,
    17'b11111101010001111,
    17'b11111101010111000,
    17'b11111101010111000,
    17'b11111101010001111,
    17'b11111101010111000,
    17'b11111101010001111,
    17'b11111101100001010,
    17'b11111101100001010,
    17'b11111101010111000,
    17'b11111101010001111,
    17'b11111101010001111,
    17'b11111101010001111,
    17'b11111101001100110,
    17'b11111101001100110,
    17'b11111101000010100,
    17'b11111101000010100,
    17'b11111101000111101,
    17'b11111101001100110,
    17'b11111101001100110,
    17'b11111101000111101,
    17'b11111101000111101,
    17'b11111101000010100,
    17'b11111101000010100,
    17'b11111101000111101,
    17'b11111101000111101,
    17'b11111101000111101,
    17'b11111101001100110,
    17'b11111101001100110,
    17'b11111101001100110,
    17'b11111101001100110,
    17'b11111101001100110,
    17'b11111101010001111,
    17'b11111101010001111,
    17'b11111101110000101,
    17'b11111110011001101,
    17'b11111110100011111,
    17'b11111110001010010,
    17'b11111110011001101,
    17'b11111111001100110,
    17'b00000000010100100,
    17'b00000001000111101,
    17'b00000000101001000,
    17'b11111110010100100,
    17'b11111011011100001,
    17'b11111000011110110,
    17'b11111001110101110,
    17'b11111010110011010,
    17'b11111011110101110,
    17'b11111100110011010,
    17'b11111101000010100,
    17'b11111100111000011,
    17'b11111101001100110,
    17'b11111100111101100,
    17'b11111101000111101,
    17'b11111101001100110,
    17'b11111101001100110,
    17'b11111101000010100,
    17'b11111101001100110,
    17'b11111101010001111,
    17'b11111101001100110,
    17'b11111101100001010,
    17'b11111101010001111,
    17'b11111101010111000,
    17'b11111101010111000,
    17'b11111101100001010,
    17'b11111101100001010,
    17'b11111101010111000,
    17'b11111101010001111,
    17'b11111101000111101,
    17'b11111101000111101,
    17'b11111101001100110,
    17'b11111101000111101,
    17'b11111101000111101,
    17'b10000000000000000,
    17'b10000000000000000,
    17'b10110000111000011,
    17'b01111100010100100,
    17'b00110111000010100,
    17'b00100010010100100,
    17'b00010010101001000,
    17'b00000100111000011,
    17'b11111110111000011,
    17'b11111011101011100,
    17'b11111010010100100,
    17'b11110111110101110,
    17'b11111000001111011,
    17'b11110100101110001,
    17'b11111010000101001,
    17'b11111110111101100,
    17'b00000111000111101,
    17'b00010100101110001,
    17'b00110010101110001,
    17'b01011000111000011,
    17'b01011011000010100,
    17'b01011001000111101,
    17'b01001011001100110,
    17'b01000000001010010,
    17'b00110110011110110,
    17'b00110000111000011,
    17'b00100111110000101,
    17'b00010101001100110,
    17'b00001100000101001,
    17'b00000000001111011,
    17'b11110001010001111,
    17'b11010110011110110,
    17'b11001101110000101,
    17'b11000111010111000,
    17'b11000011000111101,
    17'b11000001001100110,
    17'b11000010010100100,
    17'b11000110000101001,
    17'b11001011000010100,
    17'b11010010111000011,
    17'b11011010010100100,
    17'b11100010001111011,
    17'b11101110000101001,
    17'b11110101001100110,
    17'b11111010101001000,
    17'b11111110101110001,
    17'b00000001100110011,
    17'b00000011101011100,
    17'b00000101010111000,
    17'b00000110011001101,
    17'b00000100111000011,
    17'b00000000001111011,
    17'b11111010111000011,
    17'b11111001010001111,
    17'b11110111101011100,
    17'b11111000011110110,
    17'b11111011011100001,
    17'b11111101010111000,
    17'b11111101011100001,
    17'b11111100010100100,
    17'b11111011000010100,
    17'b11111010010100100,
    17'b11111011000111101,
    17'b11111110000101001,
    17'b00000000000000000,
    17'b00000001100001010,
    17'b00000010000101001,
    17'b00000010000101001,
    17'b00000001010111000,
    17'b00000001000111101,
    17'b11111111110101110,
    17'b11111101100110011,
    17'b11111100110011010,
    17'b11111100100011111,
    17'b11111100010100100,
    17'b11111101100110011,
    17'b11111100111101100,
    17'b11111100101110001,
    17'b11111110110011010,
    17'b00000000111000011,
    17'b00000000101110001,
    17'b00000000001111011,
    17'b11111111101011100,
    17'b11111111001100110,
    17'b11111110111000011,
    17'b11111110110011010,
    17'b11111110110011010,
    17'b11111111000111101,
    17'b11111111000010100,
    17'b11111110110011010,
    17'b11111110101110001,
    17'b11111110011001101,
    17'b11111110000101001,
    17'b11111101110000101,
    17'b11111101100001010,
    17'b11111101001100110,
    17'b11111101000010100,
    17'b11111101000111101,
    17'b11111110000101001,
    17'b11111110111101100,
    17'b11111110011110110,
    17'b11111110100011111,
    17'b11111110100011111,
    17'b11111110100011111,
    17'b11111111110101110,
    17'b00000010011001101,
    17'b00000011011100001,
    17'b00000100000000000,
    17'b00000011111010111,
    17'b00000011101011100,
    17'b11101001000010100,
    17'b10001010111000011,
    17'b10001100000000000,
    17'b11000000111000011,
    17'b11010001010111000,
    17'b11100001110101110,
    17'b00011011101011100,
    17'b00010101101011100,
    17'b00001110001010010,
    17'b00000110011110110,
    17'b11111011011100001,
    17'b11110001010001111,
    17'b11100111100001010,
    17'b11100111000010100,
    17'b11100110000101001,
    17'b11100100100011111,
    17'b11100011000111101,
    17'b11100101101011100,
    17'b11101101110101110,
    17'b11110101101011100,
    17'b11111001101011100,
    17'b11111101100001010,
    17'b00100111110101110,
    17'b01100010001010010,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01011110001010010,
    17'b00101000000101001,
    17'b11111100100011111,
    17'b11100011100001010,
    17'b11100000011110110,
    17'b11101111110101110,
    17'b00000101110000101,
    17'b00010111110000101,
    17'b00011110111000011,
    17'b00010111111010111,
    17'b00001111000010100,
    17'b00001011011100001,
    17'b00001111110101110,
    17'b00011001000111101,
    17'b00011010010100100,
    17'b00011101110000101,
    17'b00100011111010111,
    17'b00100111011100001,
    17'b00100110111000011,
    17'b00100011101011100,
    17'b00100000101110001,
    17'b00011111100001010,
    17'b00100000000000000,
    17'b00100001110101110,
    17'b00100100001111011,
    17'b00100011111010111,
    17'b00100101010111000,
    17'b00100111000010100,
    17'b00100101101011100,
    17'b00100011011100001,
    17'b00011111011100001,
    17'b00011000111101100,
    17'b00010101010111000,
    17'b00010001010001111,
    17'b00001110011110110,
    17'b00001100110011010,
    17'b00001010101001000,
    17'b00001001010001111,
    17'b00001001011100001,
    17'b00001011000111101,
    17'b00001100001010010,
    17'b00001100011001101,
    17'b00001011000111101,
    17'b00001010000000000,
    17'b00001001100001010,
    17'b00001001110000101,
    17'b00001011010001111,
    17'b00001100000000000,
    17'b00001110011110110,
    17'b00001110111101100,
    17'b11110010111000011,
    17'b11011000001010010,
    17'b11010101101011100,
    17'b11110010111101100,
    17'b00010001000111101,
    17'b00101101100110011,
    17'b00111111110101110,
    17'b01000011110000101,
    17'b01000011001100110,
    17'b01000110000101001,
    17'b01000101101011100,
    17'b01000000100011111,
    17'b01000010101001000,
    17'b00111101000010100,
    17'b00110011100001010,
    17'b00110001101011100,
    17'b00100000111101100,
    17'b00101010111101100,
    17'b00110101000010100,
    17'b00110101110101110,
    17'b00110011010111000,
    17'b00100100010100100,
    17'b00011010111000011,
    17'b00001110000101001,
    17'b00000101111010111,
    17'b11111011010001111,
    17'b11110111000010100,
    17'b11110101001100110,
    17'b11110100101110001,
    17'b11110010010100100,
    17'b11101111110101110,
    17'b11101110010100100,
    17'b11101001110101110,
    17'b11100010111101100,
    17'b11011110111000011,
    17'b11011101100110011,
    17'b11011010101110001,
    17'b11011100010100100,
    17'b00001011101011100,
    17'b01010111001100110,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111110010100100,
    17'b01011000010100100,
    17'b00111100001010010,
    17'b00100101100001010,
    17'b00010001001100110,
    17'b00000100011110110,
    17'b00000100010100100,
    17'b00001110001111011,
    17'b00010011110101110,
    17'b00010001000111101,
    17'b00001010101001000,
    17'b00001000011110110,
    17'b00001000101001000,
    17'b00001001101011100,
    17'b00001100100011111,
    17'b00011000100011111,
    17'b00100001010111000,
    17'b00101001000111101,
    17'b00101101000111101,
    17'b00110011000111101,
    17'b00110010111000011,
    17'b00101101110000101,
    17'b00100111010111000,
    17'b00100101000010100,
    17'b00100011101011100,
    17'b00100000100011111,
    17'b00011110011110110,
    17'b00011111000010100,
    17'b00100101010111000,
    17'b00101010000101001,
    17'b00110000000101001,
    17'b00110101101011100,
    17'b00110111100110011,
    17'b00110010100011111,
    17'b00101110011001101,
    17'b00101001101011100,
    17'b00100110111000011,
    17'b00100100110011010,
    17'b00100001110000101,
    17'b00011101110000101,
    17'b00011001010001111,
    17'b00010011101011100,
    17'b00010000101110001,
    17'b00001111111010111,
    17'b00010001001100110,
    17'b00010011010111000,
    17'b00011000100011111,
    17'b00011101110101110,
    17'b00100101001100110,
    17'b00101100101001000,
    17'b00110111111010111,
    17'b00111110011110110,
    17'b01000110011110110,
    17'b01001101110000101,
    17'b01010110000000000,
    17'b01011110011001101,
    17'b01100101011100001,
    17'b01101010101001000,
    17'b01101101011100001,
    17'b01101110000000000,
    17'b01101101011100001,
    17'b01101100110011010,
    17'b01101010111101100,
    17'b01101000110011010,
    17'b01100110010100100,
    17'b01100100101001000,
    17'b01100101010111000,
    17'b01100111101011100,
    17'b01101000010100100,
    17'b01100111100001010,
    17'b01100101110101110,
    17'b01100011100001010,
    17'b01100010001010010,
    17'b01100000110011010,
    17'b01011111100110011,
    17'b01011110001010010,
    17'b01011100011001101,
    17'b01011100000000000,
    17'b01011100000101001,
    17'b01011101010001111,
    17'b01100000011001101,
    17'b01101000001010010,
    17'b01101000010100100,
    17'b01100111100110011,
    17'b01100110001010010,
    17'b01100110011001101,
    17'b01101000000101001,
    17'b01101100101001000,
    17'b01101000101001000,
    17'b01101010000101001,
    17'b01101101101011100,
    17'b01101101010111000,
    17'b01101100100011111,
    17'b01101101011100001,
    17'b01101100111101100,
    17'b01101000111000011,
    17'b01011011001100110,
    17'b01001100111000011,
    17'b01010101010111000,
    17'b01011110011001101,
    17'b01011010110011010,
    17'b01010110011110110,
    17'b01010100010100100,
    17'b01001100100011111,
    17'b01000000111101100,
    17'b00111000111000011,
    17'b01000001101011100,
    17'b01001010000000000,
    17'b01001111110101110,
    17'b01010100001111011,
    17'b01010101001100110,
    17'b01010100001010010,
    17'b01010010011110110,
    17'b01010000101110001,
    17'b01001111011100001,
    17'b01001110000000000,
    17'b01001101110101110,
    17'b01001011110000101,
    17'b01001000111101100,
    17'b01001001010001111,
    17'b01000110101001000,
    17'b01000101110101110,
    17'b01000110000101001,
    17'b01000111000111101,
    17'b01000110101110001,
    17'b01000110011001101,
    17'b01000111110000101,
    17'b01000110101001000,
    17'b01000101010001111,
    17'b01000110110011010,
    17'b01000111110000101,
    17'b01001010011001101,
    17'b01001000000000000,
    17'b01000111010001111,
    17'b01000011001100110,
    17'b01000000100011111,
    17'b00111110101110001,
    17'b00111100000000000,
    17'b00110111010001111,
    17'b00110011100110011,
    17'b00110000010100100,
    17'b00101101000010100,
    17'b00101010111000011,
    17'b00101010101001000,
    17'b00101010010100100,
    17'b00101010000101001,
    17'b00101010011110110,
    17'b00101001100110011,
    17'b00101000001111011,
    17'b00100110101110001,
    17'b00100011011100001,
    17'b00100001010111000,
    17'b00011110001010010,
    17'b00011011111010111,
    17'b00011010011110110,
    17'b00011001101011100,
    17'b00011000100011111,
    17'b00010101100001010,
    17'b00010010100011111,
    17'b00010000010100100,
    17'b00001110000000000,
    17'b00001001100001010,
    17'b00000101100001010,
    17'b00000001110101110,
    17'b11111110110011010,
    17'b11111100001111011,
    17'b11111010001010010,
    17'b11111000111101100,
    17'b11111000010100100,
    17'b11110111011100001,
    17'b11110101100001010,
    17'b11110011100110011,
    17'b11110000111101100,
    17'b11101101110101110,
    17'b11101001110000101,
    17'b11100111000111101,
    17'b11100101010111000,
    17'b11100100000000000,
    17'b11100001101011100,
    17'b11100000111000011,
    17'b11011011111010111,
    17'b11010110101001000,
    17'b11010011100110011,
    17'b11001101101011100,
    17'b11001000110011010,
    17'b11000110000000000,
    17'b11000000011110110,
    17'b10111100000101001,
    17'b10111000111101100,
    17'b10110110000000000,
    17'b10110011101011100,
    17'b10110001110000101,
    17'b10101111001100110,
    17'b10101101111010111,
    17'b10101100101001000,
    17'b10101100001010010,
    17'b10101011010111000,
    17'b10101011100001010,
    17'b10101011100001010,
    17'b10101100010100100,
    17'b10101100101110001,
    17'b10101101100110011,
    17'b10101110011110110,
    17'b10101110101001000,
    17'b10101110110011010,
    17'b10101110010100100,
    17'b10101101110101110,
    17'b10101101111010111,
    17'b10101101010111000,
    17'b10101101000111101,
    17'b10101100011110110,
    17'b10101100000000000,
    17'b10101011101011100,
    17'b10101011110000101,
    17'b10101100000000000,
    17'b10101100101001000,
    17'b10101101010111000,
    17'b10101110000000000,
    17'b10101111000111101,
    17'b10101111010001111,
    17'b10101111100001010,
    17'b10101110111000011,
    17'b10101101010001111,
    17'b10101011101011100,
    17'b10101001110101110,
    17'b10100111111010111,
    17'b10100110101110001,
    17'b10100100101001000,
    17'b10100011010111000,
    17'b10100010100011111,
    17'b10100001111010111,
    17'b10100001011100001,
    17'b10100001011100001,
    17'b10100010001111011,
    17'b10100010111101100,
    17'b10100100000000000,
    17'b10100101110000101,
    17'b10100111010111000,
    17'b10101001010001111,
    17'b10101011011100001,
    17'b10101111000111101,
    17'b10110010011110110,
    17'b10110100111000011,
    17'b10110110111101100,
    17'b10111011011100001,
    17'b10111100001111011,
    17'b10111001000111101,
    17'b10111000001010010,
    17'b10111001000111101,
    17'b10111001100110011,
    17'b10110110111101100,
    17'b10110110000101001,
    17'b10110111000111101,
    17'b10110101111010111,
    17'b10110111000111101,
    17'b10110110011001101,
    17'b10110101111010111,
    17'b10111000111000011,
    17'b10111011110101110,
    17'b10111110111101100,
    17'b11000010001111011,
    17'b11000100100011111,
    17'b11000110101110001,
    17'b11001010001111011,
    17'b11001110001010010,
    17'b11010100010100100,
    17'b11011001100001010,
    17'b11100010101110001,
    17'b11110001010111000,
    17'b11111101001100110,
    17'b00000000111101100,
    17'b00000011001100110,
    17'b00001000100011111,
    17'b00011101100001010,
    17'b00101111010111000,
    17'b00111011011100001,
    17'b00110100110011010,
    17'b00000010001010010,
    17'b11011100111000011,
    17'b11011010111000011,
    17'b11101101110000101,
    17'b00001111100001010,
    17'b01111111111111111,
    17'b01010000010100100,
    17'b00010011101011100,
    17'b00000010001111011,
    17'b00000010001010010,
    17'b11110100001010010,
    17'b11011101110000101,
    17'b11011000111000011,
    17'b11100000000101001,
    17'b11101110001010010,
    17'b11110111001100110,
    17'b11111100110011010,
    17'b00000000011001101,
    17'b11110110001111011,
    17'b11110011111010111,
    17'b11110100000000000,
    17'b11110101110101110,
    17'b11111100011001101,
    17'b11110100011110110,
    17'b11110010001010010,
    17'b11111000011001101,
    17'b00001011000010100,
    17'b00011110000101001,
    17'b00100100101001000,
    17'b00011011100110011,
    17'b00010011000010100,
    17'b00001110010100100,
    17'b00000100111000011,
    17'b11111011111010111,
    17'b11101010111101100,
    17'b11011000110011010,
    17'b11001111000111101,
    17'b11001000000101001,
    17'b11001010110011010,
    17'b11010001110101110,
    17'b11010000101110001,
    17'b11010000001111011,
    17'b11011101011100001,
    17'b11100101111010111,
    17'b11110100001111011,
    17'b00000111111010111,
    17'b00000111110101110,
    17'b11110011111010111,
    17'b11100111000010100,
    17'b11110010101110001,
    17'b11110110001010010,
    17'b11110001101011100,
    17'b11101110000000000,
    17'b11101010001111011,
    17'b11101011101011100,
    17'b11110000101110001,
    17'b11101111011100001,
    17'b11101000101001000,
    17'b11100010100011111,
    17'b11011011010111000,
    17'b11011010111000011,
    17'b11011001110000101,
    17'b11100001000111101,
    17'b11011111000010100,
    17'b11100000111101100,
    17'b11010111000111101,
    17'b11011111011100001,
    17'b11100101111010111,
    17'b11101101111010111,
    17'b11111000001111011,
    17'b11111010100011111,
    17'b11111001001100110,
    17'b11110010110011010,
    17'b11101011100110011,
    17'b11101011100001010,
    17'b11101110000000000,
    17'b11110000010100100,
    17'b11101110001111011,
    17'b11101101010001111,
    17'b11110000110011010,
    17'b11110111000010100,
    17'b11110111101011100,
    17'b11110010011001101,
    17'b11101101010001111,
    17'b11101000001010010,
    17'b11100010101110001,
    17'b11011101010111000,
    17'b11011000000000000,
    17'b11010001100001010,
    17'b11001110000000000,
    17'b11001011001100110,
    17'b11001001100001010,
    17'b11001001110000101,
    17'b11001011100110011,
    17'b11001110011001101,
    17'b11010001001100110,
    17'b11010101010001111,
    17'b11011001011100001,
    17'b11011101000111101,
    17'b11100000011110110,
    17'b11100100001111011,
    17'b11100110101110001,
    17'b11101000010100100,
    17'b11101001101011100,
    17'b11101100011110110,
    17'b11101100101001000,
    17'b11101110101110001,
    17'b11101111111010111,
    17'b11110001010001111,
    17'b11110011100001010,
    17'b11110110101110001,
    17'b11111100110011010,
    17'b00000010001111011,
    17'b00001000010100100,
    17'b00000111111010111,
    17'b00001001010111000,
    17'b00001010000000000,
    17'b00001010000101001,
    17'b00001001000111101,
    17'b00000110011001101,
    17'b00000011111010111,
    17'b00000011101011100,
    17'b00000100001010010,
    17'b11111101110000101,
    17'b00000000011001101,
    17'b11111111110101110,
    17'b11111100000101001,
    17'b00000001110000101,
    17'b11111111000111101,
    17'b11111100000000000,
    17'b11110011111010111,
    17'b11111011101011100,
    17'b11101100011001101,
    17'b11100111011100001,
    17'b11011110111101100,
    17'b11011110101110001,
    17'b11001111010111000,
    17'b11011010101110001,
    17'b11010100111000011,
    17'b11001110011110110,
    17'b11010010101110001,
    17'b11001110011110110,
    17'b11001011110000101,
    17'b11000101001100110,
    17'b11001110100011111,
    17'b11001110011110110,
    17'b11001011101011100,
    17'b11001101000010100,
    17'b11001011100110011,
    17'b11001000111000011,
    17'b11001001111010111,
    17'b11001101100110011,
    17'b11010010000101001,
    17'b11010101111010111,
    17'b11010110111000011,
    17'b11010111111010111,
    17'b11011001011100001,
    17'b11011001010111000,
    17'b11011111010111000,
    17'b11100001110000101,
    17'b11100101000010100,
    17'b11100111111010111,
    17'b11100001010001111,
    17'b11011111001100110,
    17'b11011110000101001,
    17'b11011100110011010,
    17'b11011010001010010,
    17'b11011010100011111,
    17'b11011010001010010,
    17'b11011001110000101,
    17'b11010111011100001,
    17'b11010101101011100,
    17'b11010111100110011,
    17'b11011000000101001,
    17'b11011000001111011,
    17'b11011001110101110,
    17'b11011000100011111,
    17'b11011001110101110,
    17'b11011000101110001,
    17'b11010110111101100,
    17'b11010110101110001,
    17'b11100010001111011,
    17'b11110010101110001,
    17'b11110011010111000,
    17'b11110000010100100,
    17'b11111000101001000,
    17'b00000000101001000,
    17'b11111110001010010,
    17'b11110101111010111,
    17'b11101110000000000,
    17'b11101010001010010,
    17'b11101000100011111,
    17'b11100011010001111,
    17'b11010100001010010,
    17'b11011110011110110,
    17'b11011101010111000,
    17'b11100101001100110,
    17'b11111000110011010,
    17'b00000011110101110,
    17'b11110001111010111,
    17'b11101010111000011,
    17'b11101101111010111,
    17'b00000110000000000,
    17'b00000011000111101,
    17'b11111000011110110,
    17'b11101111001100110,
    17'b11011011100110011,
    17'b10111110010100100,
    17'b10110111100110011,
    17'b11100110000101001,
    17'b11101101001100110,
    17'b00001010000101001,
    17'b00100001111010111,
    17'b00101000101001000,
    17'b00011011000111101,
    17'b00000111010111000,
    17'b00000011110000101,
    17'b00000100000101001,
    17'b00000100100011111,
    17'b00000010011001101,
    17'b00000001000010100,
    17'b11111110000000000,
    17'b11111011011100001,
    17'b11111011111010111,
    17'b11111011110000101,
    17'b11111010100011111,
    17'b11110111011100001,
    17'b11110101100110011,
    17'b11110110000000000,
    17'b11110010011001101,
    17'b11100101010111000,
    17'b11010111111010111,
    17'b10111111110101110,
    17'b11000111011100001,
    17'b11011111010111000,
    17'b11110111110101110,
    17'b00010000111101100,
    17'b00011011010001111,
    17'b00011100001010010,
    17'b00010010101001000,
    17'b00000011100001010,
    17'b11110111101011100,
    17'b11110001100001010,
    17'b11101110100011111,
    17'b11101110101001000,
    17'b11101110011110110,
    17'b11110100001010010,
    17'b11111100010100100,
    17'b00000100000101001,
    17'b00000101000010100,
    17'b00000101000111101,
    17'b00000111100001010,
    17'b00000111101011100,
    17'b00000011001100110,
    17'b11111101000111101,
    17'b11111001110101110,
    17'b11110101010111000,
    17'b11110100000101001,
    17'b11110000011110110,
    17'b11101010010100100,
    17'b11011100001010010,
    17'b11000011111010111,
    17'b11000000010100100,
    17'b11010101011100001,
    17'b11011111100110011,
    17'b11101011011100001,
    17'b11111101011100001,
    17'b00000000011110110,
    17'b11111100111000011,
    17'b11111010100011111,
    17'b11110110000000000,
    17'b11110010011001101,
    17'b11110000110011010,
    17'b11101110100011111,
    17'b11101011100001010,
    17'b11100111111010111,
    17'b11100100110011010,
    17'b11100011000010100,
    17'b11100001111010111,
    17'b11100001100110011,
    17'b11100001111010111,
    17'b11100001011100001,
    17'b11100010010100100,
    17'b11101000000101001,
    17'b00000000111101100,
    17'b00100001110101110,
    17'b00011010010100100,
    17'b00001001111010111,
    17'b11111001010111000,
    17'b11100010111101100,
    17'b11011011010001111,
    17'b11011001010111000,
    17'b11011100110011010,
    17'b11001111100001010,
    17'b11000011100110011,
    17'b10111110101110001,
    17'b11000011001100110,
    17'b11011001010111000,
    17'b11100101110101110,
    17'b11101001101011100,
    17'b11101010000000000,
    17'b11101110111000011,
    17'b11110010011001101,
    17'b11110001110101110,
    17'b11101111110101110,
    17'b11101111011100001,
    17'b11101111110101110,
    17'b11101111101011100,
    17'b11101101100001010,
    17'b11101100100011111,
    17'b11110010101001000,
    17'b11110101001100110,
    17'b11110101011100001,
    17'b11110111101011100,
    17'b11111011000010100,
    17'b11111110011001101,
    17'b00000000110011010,
    17'b00000011000111101,
    17'b00000100011110110,
    17'b00000101010111000,
    17'b00000101111010111,
    17'b00000110101110001,
    17'b00001000100011111,
    17'b00001001111010111,
    17'b00001010101110001,
    17'b00001011000010100,
    17'b00001011010111000,
    17'b00001011000111101,
    17'b00001010010100100,
    17'b00001001000111101,
    17'b00000111011100001,
    17'b00000110111101100,
    17'b00000111000010100,
    17'b00000110111101100,
    17'b00000101110101110,
    17'b00000011001100110,
    17'b00000000100011111,
    17'b11111110011001101,
    17'b11111100110011010,
    17'b11111011011100001,
    17'b11111011010001111,
    17'b11111010111101100,
    17'b11111011001100110,
    17'b11111011110101110,
    17'b11111100111000011,
    17'b11111110011001101,
    17'b00000001000010100,
    17'b00000100011001101,
    17'b00001000111000011,
    17'b00001100001010010,
    17'b00001110101001000,
    17'b00010000001010010,
    17'b00010001000010100,
    17'b00010000100011111,
    17'b00001100011001101,
    17'b00001010111101100,
    17'b00001101110000101,
    17'b00001110011110110,
    17'b00001110110011010,
    17'b00001011010001111,
    17'b00001010111000011,
    17'b00001010111101100,
    17'b00001010111101100,
    17'b00001010110011010,
    17'b00001001101011100,
    17'b00000111010111000,
    17'b00000100011001101,
    17'b11111111110101110,
    17'b11111101001100110,
    17'b11111011001100110,
    17'b11111010000101001,
    17'b11111001111010111,
    17'b11111011100001010,
    17'b00000001110000101,
    17'b00001001100001010,
    17'b00010001010111000,
    17'b00010101011100001,
    17'b00011000000101001,
    17'b00011001100110011,
    17'b00011011010001111,
    17'b00011101000010100,
    17'b00100010011001101,
    17'b00101100001010010,
    17'b00111000001111011,
    17'b00111101010001111,
    17'b00111100111000011,
    17'b00111000001111011,
    17'b00110011000010100,
    17'b00101110111000011,
    17'b00101110101001000,
    17'b00110000011001101,
    17'b00110010001010010,
    17'b00110011010001111,
    17'b00110100100011111,
    17'b00110101100001010,
    17'b00110110111101100,
    17'b00110111011100001,
    17'b00110110000000000,
    17'b00110011000010100,
    17'b00101110101110001,
    17'b00101010111101100,
    17'b00100111001100110,
    17'b00100100111000011,
    17'b00100100011110110,
    17'b00100101001100110,
    17'b00100110001010010,
    17'b00100111010001111,
    17'b00100111110101110,
    17'b00100111111010111,
    17'b00100110011110110,
    17'b00100100100011111,
    17'b00100010011001101,
    17'b00100000000101001,
    17'b00011111101011100,
    17'b00011111110000101,
    17'b00100000001010010,
    17'b00100000110011010,
    17'b00100010010100100,
    17'b00100011010001111,
    17'b00100100101001000,
    17'b00100101100110011,
    17'b00100110000000000,
    17'b00100101100110011,
    17'b00100100100011111,
    17'b00100011001100110,
    17'b00100001010001111,
    17'b00011111011100001,
    17'b00011110111101100,
    17'b00011111010001111,
    17'b00100000000101001,
    17'b00100001110101110,
    17'b00100010100011111,
    17'b00100010001010010,
    17'b00100000110011010,
    17'b00100001010001111,
    17'b00011111010001111,
    17'b00011110011001101,
    17'b00011111100001010,
    17'b00011111100110011,
    17'b00011011100110011,
    17'b00010111110000101,
    17'b00010101010111000,
    17'b00010010101001000,
    17'b00010010000101001,
    17'b00010001111010111,
    17'b00010001010111000,
    17'b00010000100011111,
    17'b00010000110011010,
    17'b00010011011100001,
    17'b00010011011100001,
    17'b00010110001010010,
    17'b00010111000010100,
    17'b00010101011100001,
    17'b00010011110101110,
    17'b00010010100011111,
    17'b00010000001111011,
    17'b00001101110000101,
    17'b00001011000111101,
    17'b00001001100001010,
    17'b00001000000101001,
    17'b00001000001010010,
    17'b00001000111000011,
    17'b00000010011110110,
    17'b00000110111000011,
    17'b00001110001111011,
    17'b00010100100011111,
    17'b00010100101110001,
    17'b00001110110011010,
    17'b11111111101011100,
    17'b11111101111010111,
    17'b00000011010001111,
    17'b00000011110101110,
    17'b11111110111000011,
    17'b11111001110101110,
    17'b11110111011100001,
    17'b11111100001010010,
    17'b00000110010100100,
    17'b00001001100110011,
    17'b00001000110011010,
    17'b00000111010001111,
    17'b00000101011100001,
    17'b00000010111000011,
    17'b00000001110000101,
    17'b00000000001111011,
    17'b11111111001100110,
    17'b11111110001111011,
    17'b11111110001111011,
    17'b11111111010001111,
    17'b00000000001111011,
    17'b00000000011001101,
    17'b11111111110000101,
    17'b11111111100110011,
    17'b11111111110101110,
    17'b11111100110011010,
    17'b11111001101011100,
    17'b11110011000010100,
    17'b11110000011001101,
    17'b11111000000000000,
    17'b11111110001111011,
    17'b11111000111000011,
    17'b11110011001100110,
    17'b11101100111101100,
    17'b11110000000000000,
    17'b11110110011110110,
    17'b00000101100110011,
    17'b00010110011001101,
    17'b00011111010001111,
    17'b00100010111000011,
    17'b00011110101001000,
    17'b00010010000101001,
    17'b00001000000000000,
    17'b11111001111010111,
    17'b11101111110101110,
    17'b11101010010100100,
    17'b11101010101110001,
    17'b11110001111010111,
    17'b11111100000000000,
    17'b00000101000010100,
    17'b00001010000101001,
    17'b00001010001111011,
    17'b00000111110101110,
    17'b00000100111101100,
    17'b00000100000101001,
    17'b00000011110000101,
    17'b00000100000101001,
    17'b00000100101110001,
    17'b00000101100110011,
    17'b00000110000101001,
    17'b00000101111010111,
    17'b00000100111000011,
    17'b00000100000101001,
    17'b00000011010111000,
    17'b00000011000010100,
    17'b00000011000111101,
    17'b00000100001010010,
    17'b00000101101011100,
    17'b00000111010001111,
    17'b00001000000101001,
    17'b00001000011110110,
    17'b00000111100001010,
    17'b00000100101110001,
    17'b00000001000010100,
    17'b11111110110011010,
    17'b11111110100011111,
    17'b11111111000111101,
    17'b11111111000111101,
    17'b11111110101001000,
    17'b11111101110000101,
    17'b11111101000111101,
    17'b11111101001100110,
    17'b11111101100110011,
    17'b11111110001010010,
    17'b11111101100001010,
    17'b11111100100011111,
    17'b11111010111101100,
    17'b11111001000010100,
    17'b11110111101011100,
    17'b11111000001010010,
    17'b11111001101011100,
    17'b00000001001100110,
    17'b00001101000010100,
    17'b00011000010100100,
    17'b00011100001010010,
    17'b00011010000101001,
    17'b00010111001100110,
    17'b00010110001111011,
    17'b00001110110011010,
    17'b00000111111010111,
    17'b00000011011100001,
    17'b00000001000010100,
    17'b11111111011100001,
    17'b11111110111101100,
    17'b11111101100001010,
    17'b11111101111010111,
    17'b11111111000111101,
    17'b00000000110011010,
    17'b00000010101001000,
    17'b00000101100110011,
    17'b00001000000101001,
    17'b00001010100011111,
    17'b00001100110011010,
    17'b00001110101001000,
    17'b00001111110101110,
    17'b00010000101001000,
    17'b00010001100001010,
    17'b00010001101011100,
    17'b00010001100110011,
    17'b00010001101011100,
    17'b00010001100001010,
    17'b00010000100011111,
    17'b00001110111101100,
    17'b00001100000000000,
    17'b00001011000010100,
    17'b00001001110101110,
    17'b00001001010001111,
    17'b00001010101001000,
    17'b00001110101110001,
    17'b00010010000101001,
    17'b00010101010001111,
    17'b00011000000000000,
    17'b00011001101011100,
    17'b00011001110000101,
    17'b00011000000101001,
    17'b00010101000010100,
    17'b00010001011100001,
    17'b00001101110000101,
    17'b00001001111010111,
    17'b00001000001010010,
    17'b00000111011100001,
    17'b00000110111101100,
    17'b00000110111000011,
    17'b00000111001100110,
    17'b00000111110101110,
    17'b00001000011110110,
    17'b00001001100001010,
    17'b00001100100011111,
    17'b00010001000111101,
    17'b00010011110000101,
    17'b00010100000101001,
    17'b00010100000000000,
    17'b00010011010001111,
    17'b00010010000000000,
    17'b00010001111010111,
    17'b00010001101011100,
    17'b00010000001111011,
    17'b00001110111101100,
    17'b00001110110011010,
    17'b00001110011001101,
    17'b00001100111000011,
    17'b00001010101001000,
    17'b00001000111000011,
    17'b00010010001111011,
    17'b00011101010001111,
    17'b00100101000111101,
    17'b00100111010111000,
    17'b00100010111000011,
    17'b00011101001100110,
    17'b00011000001010010,
    17'b00010011100001010,
    17'b00010010010100100,
    17'b00010100111000011,
    17'b00010111011100001,
    17'b00011000101110001,
    17'b00011010001010010,
    17'b00011011000010100,
    17'b00011011010001111,
    17'b00011011101011100,
    17'b00011100111101100,
    17'b00011110001010010,
    17'b00011110011110110,
    17'b00011100010100100,
    17'b00100011000010100,
    17'b00101001100001010,
    17'b00100101101011100,
    17'b00100001000010100,
    17'b00011111111010111,
    17'b00011111001100110,
    17'b00011110111101100,
    17'b00100000111000011,
    17'b00100011110000101,
    17'b00100110100011111,
    17'b00100111111010111,
    17'b00101001000111101,
    17'b00101110100011111,
    17'b00101111000111101,
    17'b00110011110000101,
    17'b00110100110011010,
    17'b00110011100110011,
    17'b00110110001010010,
    17'b00110110110011010,
    17'b00110010111000011,
    17'b00101001110101110,
    17'b00011110101110001,
    17'b00010101110000101,
    17'b00001110101001000,
    17'b00001100100011111,
    17'b00001100011001101,
    17'b00001110001111011,
    17'b00010011011100001,
    17'b00010111010001111,
    17'b00011001100001010,
    17'b00011001011100001,
    17'b00010100011001101,
    17'b00010100000000000,
    17'b00010010111101100,
    17'b00001110110011010,
    17'b00001010111000011,
    17'b00001010100011111,
    17'b00001010110011010,
    17'b00001011010001111,
    17'b00001011110101110,
    17'b00001100110011010,
    17'b00001101100110011,
    17'b00001110101001000,
    17'b00010000000000000,
    17'b00010010000000000,
    17'b00010011000010100,
    17'b00010010111101100,
    17'b00010010000000000,
    17'b00010000101110001,
    17'b00001110000101001,
    17'b00001011011100001,
    17'b00001000001111011,
    17'b00000101000010100,
    17'b00000010000000000,
    17'b00000001000010100,
    17'b00000000100011111,
    17'b00000000111101100,
    17'b00000010001111011,
    17'b00000101010111000,
    17'b00001000101001000,
    17'b00001011110000101,
    17'b00001101100110011,
    17'b00001110011001101,
    17'b00001110101110001,
    17'b00001101010111000,
    17'b00001000011110110,
    17'b00000001010111000,
    17'b11111010001111011,
    17'b11110101101011100,
    17'b11110111000111101,
    17'b11111011011100001,
    17'b00000000100011111,
    17'b00000101010001111,
    17'b00001010100011111,
    17'b00001110111000011,
    17'b00010100000000000,
    17'b00011000111101100,
    17'b00011100101110001,
    17'b00011101011100001,
    17'b00011101010001111,
    17'b00011100111000011,
    17'b00011101110000101,
    17'b00011111101011100,
    17'b00100000100011111,
    17'b00100001001100110,
    17'b00100101000111101,
    17'b00100111000010100,
    17'b00100101010001111,
    17'b00100111010001111,
    17'b00100010011001101,
    17'b00011010101110001,
    17'b00010101010111000,
    17'b00011101010111000,
    17'b00100010101110001,
    17'b00100101101011100,
    17'b00100110110011010,
    17'b00101001100001010,
    17'b00101001100110011,
    17'b00100111100001010,
    17'b00100111000010100,
    17'b00101000011110110,
    17'b00101010101110001,
    17'b00101000101110001,
    17'b00101101000111101,
    17'b00110010011001101,
    17'b00110101000111101,
    17'b00111010111101100,
    17'b01000010001111011,
    17'b01001011011100001,
    17'b01001011110000101,
    17'b01001011000111101,
    17'b01001001011100001,
    17'b01001000000000000,
    17'b01000111001100110,
    17'b01000100101001000,
    17'b01000011010001111,
    17'b01000101000010100,
    17'b01000111100001010,
    17'b01001010010100100,
    17'b01001101001100110,
    17'b01010000000101001,
    17'b01010010011001101,
    17'b01010010100011111,
    17'b01010000100011111,
    17'b01001101011100001,
    17'b01001010101001000,
    17'b01000111110101110,
    17'b01000101100110011,
    17'b01000100010100100,
    17'b01000100110011010,
    17'b01001001010001111,
    17'b01001111011100001,
    17'b01010011111010111,
    17'b01011010100011111,
    17'b01011111010111000,
    17'b01011111000111101,
    17'b01011110110011010,
    17'b01010111100110011,
    17'b01010011011100001,
    17'b01010001010111000,
    17'b01010001011100001,
    17'b01010011100110011,
    17'b01010100011001101,
    17'b01010100101001000,
    17'b01010110000101001,
    17'b01011000101001000,
    17'b01011010000000000,
    17'b01011011000010100,
    17'b01011011110101110,
    17'b01011011111010111,
    17'b01011010111000011,
    17'b01011001010001111,
    17'b01011000000101001,
    17'b01011000001111011,
    17'b01100000000101001,
    17'b01011000111101100,
    17'b01000101000010100,
    17'b01001001000010100,
    17'b01001000100011111,
    17'b01000101011100001,
    17'b01000001000111101,
    17'b00111111100110011,
    17'b00111001001100110,
    17'b00110110101110001,
    17'b00110111110000101,
    17'b00110110111000011,
    17'b00111011000111101,
    17'b00111010011110110,
    17'b00110111101011100,
    17'b00111010100011111,
    17'b00111001000111101,
    17'b00111000001010010,
    17'b00111000000101001,
    17'b00110110111000011,
    17'b00110101100001010,
    17'b00110111101011100,
    17'b00111001111010111,
    17'b00111010010100100,
    17'b00111010000101001,
    17'b00110101100001010,
    17'b00101011110101110,
    17'b00011100001111011,
    17'b00010001100001010,
    17'b00001111111010111,
    17'b00001010100011111,
    17'b00001110001111011,
    17'b00010000101001000,
    17'b00011010001111011,
    17'b00110000011001101,
    17'b00111000001010010,
    17'b00101110000000000,
    17'b00011001110101110,
    17'b00001001010001111,
    17'b11111101000010100,
    17'b11111000101110001,
    17'b11110100101110001,
    17'b11110000001010010,
    17'b11101101110000101,
    17'b11110000000000000,
    17'b11110010011110110,
    17'b11110100001111011,
    17'b11110011000111101,
    17'b11101100101110001,
    17'b11100110110011010,
    17'b11101011111010111,
    17'b11101101010111000,
    17'b11101111000010100,
    17'b11110000011110110,
    17'b11110000101001000,
    17'b11110000000000000,
    17'b11101111000010100,
    17'b11101110000101001,
    17'b11101100111101100,
    17'b11101100011110110,
    17'b11101100000101001,
    17'b11101011111010111,
    17'b11101100101110001,
    17'b11101101100110011,
    17'b11101110010100100,
    17'b11101111010001111,
    17'b11110000111000011,
    17'b11110010110011010,
    17'b11110100110011010,
    17'b11110101101011100,
    17'b11110100111101100,
    17'b11110101100110011,
    17'b11110101110101110,
    17'b11110110000000000,
    17'b11111001001100110,
    17'b00000001100001010,
    17'b00001001011100001,
    17'b00000110100011111,
    17'b11111110000101001,
    17'b11111001011100001,
    17'b11110011010111000,
    17'b11101100000000000,
    17'b11101001111010111,
    17'b11101001010111000,
    17'b11101000110011010,
    17'b11100010101001000,
    17'b11011001011100001,
    17'b11010001010001111,
    17'b11001010001010010,
    17'b11000100000101001,
    17'b10111110111000011,
    17'b10111101111010111,
    17'b11000011111010111,
    17'b11001011110101110,
    17'b11010100000000000,
    17'b11011011000111101,
    17'b11100011000010100,
    17'b11101000011001101,
    17'b11101101001100110,
    17'b11110000111101100,
    17'b11110011000010100,
    17'b11110010011001101,
    17'b11110000101001000,
    17'b11101111100110011,
    17'b11110000011110110,
    17'b11110010100011111,
    17'b11110101010001111,
    17'b11111001001100110,
    17'b11111100010100100,
    17'b11111111000010100,
    17'b00000000010100100,
    17'b00000011001100110,
    17'b00000110010100100,
    17'b00000111100110011,
    17'b00000111010001111,
    17'b00000101100110011,
    17'b11111101000010100,
    17'b11111100000000000,
    17'b11111010111101100,
    17'b11111010000101001,
    17'b11110111110101110,
    17'b11110011100110011,
    17'b11101101010111000,
    17'b11101001100110011,
    17'b11100111000111101,
    17'b11100111100001010,
    17'b11101010110011010,
    17'b11101101101011100,
    17'b11110000000000000,
    17'b11110010011001101,
    17'b11110100000101001,
    17'b11110110101001000,
    17'b11111010000101001,
    17'b11111110111101100,
    17'b00000001111010111,
    17'b00000011011100001,
    17'b00000011010111000,
    17'b00000010000000000,
    17'b00000000111000011,
    17'b00000001011100001,
    17'b00000010111101100,
    17'b00000100101001000,
    17'b00000110101110001,
    17'b00000111010111000,
    17'b00000110011110110,
    17'b00000100001111011,
    17'b00000000111000011,
    17'b00000000000101001,
    17'b00000000100011111,
    17'b00000000111101100,
    17'b00000000001111011,
    17'b11111111010001111,
    17'b11111110100011111,
    17'b11111101000010100,
    17'b11111010111000011,
    17'b11111011010001111,
    17'b11111101100001010,
    17'b11111111011100001,
    17'b11111111001100110,
    17'b11111110101001000,
    17'b11111110000000000,
    17'b11111101100001010,
    17'b11111101010001111,
    17'b11111110000000000,
    17'b11111111010111000,
    17'b00000001000111101,
    17'b00000001111010111,
    17'b00000010111000011,
    17'b00000011111010111,
    17'b00000100011001101,
    17'b00000011110000101,
    17'b00000011010111000,
    17'b00000010110011010,
    17'b00000001110000101,
    17'b00000001001100110,
    17'b00000001010111000,
    17'b00000010001010010,
    17'b00000010111000011,
    17'b00000011100001010,
    17'b00000011011100001,
    17'b00000011001100110,
    17'b00000011001100110,
    17'b00000011000010100,
    17'b00000010101110001,
    17'b00000010001111011,
    17'b00000001110000101,
    17'b00000000110011010,
    17'b11111111010111000,
    17'b11111101100110011,
    17'b11111100001010010,
    17'b11111011110000101,
    17'b11111100110011010,
    17'b11111101011100001,
    17'b11111111010111000,
    17'b00000001111010111,
    17'b00000001111010111,
    17'b11111110111000011,
    17'b11111100101001000,
    17'b11111011010001111,
    17'b11111001001100110,
    17'b11110101100001010,
    17'b11110011001100110,
    17'b11110001111010111,
    17'b11110001000010100,
    17'b11101111010111000,
    17'b11110000001010010,
    17'b11110001001100110,
    17'b11110010000101001,
    17'b11110010111000011,
    17'b11110011010001111,
    17'b11110101110000101,
    17'b11110110010100100,
    17'b11110110101001000,
    17'b11110110000101001,
    17'b11110110011110110,
    17'b11111000111101100,
    17'b11111001011100001,
    17'b11111010000101001,
    17'b11111011001100110,
    17'b11111110001111011,
    17'b11111110101001000,
    17'b11111110011110110,
    17'b00000110101001000,
    17'b00001011100110011,
    17'b00010000011110110,
    17'b00011100000101001,
    17'b00101100001010010,
    17'b01001101010111000,
    17'b01011000001111011,
    17'b01000110001010010,
    17'b00101100111000011,
    17'b00010110011110110,
    17'b00000101110101110,
    17'b11111100110011010,
    17'b11110101111010111,
    17'b11101011110101110,
    17'b11100010011110110,
    17'b11011101000010100,
    17'b11011110000000000,
    17'b11100010110011010,
    17'b11100001110101110,
    17'b11101100001111011,
    17'b11110101111010111,
    17'b11110111010111000,
    17'b11110110000101001,
    17'b11110101010001111,
    17'b11110110001010010,
    17'b11111010000101001,
    17'b11111101010001111,
    17'b11111111011100001,
    17'b00000001010001111,
    17'b00000010101110001,
    17'b00000100000101001,
    17'b00000000001111011,
    17'b11111101110000101,
    17'b00000110011110110,
    17'b00000010001010010,
    17'b11110000001010010,
    17'b11101000110011010,
    17'b11100101010001111,
    17'b11100011011100001,
    17'b11100110010100100,
    17'b11101001000010100,
    17'b11100111011100001,
    17'b11100010101001000,
    17'b11011110111000011,
    17'b11011100101110001,
    17'b11100001000111101,
    17'b11101101100001010,
    17'b11110011011100001,
    17'b11110011000010100,
    17'b11110100000101001,
    17'b11110100111101100,
    17'b11110011110101110,
    17'b11110010001111011,
    17'b11101110101001000,
    17'b11101101010111000,
    17'b11110000011110110,
    17'b11101101101011100,
    17'b11110000000000000,
    17'b11110111010111000,
    17'b00000001000010100,
    17'b00000011100001010,
    17'b00000010001010010,
    17'b00000000000101001,
    17'b11111110001010010,
    17'b11111011010001111,
    17'b11110111100001010,
    17'b11110110011110110,
    17'b11110000100011111,
    17'b11101011010001111,
    17'b11100100110011010,
    17'b11100101010001111,
    17'b11100110011110110,
    17'b11101001100001010,
    17'b11111000111000011,
    17'b00001101011100001,
    17'b00001000111101100,
    17'b00000011110000101,
    17'b00000000001010010,
    17'b11111100111101100,
    17'b11111010011110110,
    17'b11111011111010111,
    17'b11111101110101110,
    17'b00000000011110110,
    17'b00000010011001101,
    17'b00000100101001000,
    17'b00000111111010111,
    17'b00001010000101001,
    17'b00001100000101001,
    17'b00001101101011100,
    17'b00001111100001010,
    17'b00010000100011111,
    17'b00010001011100001,
    17'b00010010011110110,
    17'b00010100100011111,
    17'b00010111000010100,
    17'b00011001110000101,
    17'b00011100101110001,
    17'b00100000011001101,
    17'b00100010010100100,
    17'b00100011001100110,
    17'b00100011011100001,
    17'b00100011100001010,
    17'b00100011100001010,
    17'b00100011100001010,
    17'b00100011000111101,
    17'b00100010100011111,
    17'b00100010001010010,
    17'b00100011111010111,
    17'b00100100110011010,
    17'b00100100100011111,
    17'b00100011101011100,
    17'b00100010011110110,
    17'b00100001100110011,
    17'b00100010001010010,
    17'b00100010111000011,
    17'b00100011000010100,
    17'b00100010110011010,
    17'b00100001010001111,
    17'b00100001101011100,
    17'b00100010001111011,
    17'b00100010000000000,
    17'b00100010011001101,
    17'b00100100001010010,
    17'b00100110101110001,
    17'b00101010000101001,
    17'b00101100100011111,
    17'b00110000000000000,
    17'b00110010101001000,
    17'b00110100110011010,
    17'b00110100110011010,
    17'b00110100001111011,
    17'b00110100011110110,
    17'b00110100000101001,
    17'b00110010111000011,
    17'b00110001111010111,
    17'b00110001010111000,
    17'b00110010101110001,
    17'b00110101110101110,
    17'b00111010110011010,
    17'b01000000100011111,
    17'b01000011100001010,
    17'b01000100001111011,
    17'b01000100001111011,
    17'b01010011100001010,
    17'b01010111100110011,
    17'b01011101000010100,
    17'b01100010011110110,
    17'b01101001011100001,
    17'b01100100011001101,
    17'b01011010111000011,
    17'b01010010111101100,
    17'b01001111001100110,
    17'b01001110101110001,
    17'b01001101010001111,
    17'b01001101011100001,
    17'b01001100000000000,
    17'b01000100001010010,
    17'b00111010110011010,
    17'b00111010100011111,
    17'b00111111100001010,
    17'b01000101010111000,
    17'b01000111100110011,
    17'b01001010000000000,
    17'b01001011110000101,
    17'b01001010110011010,
    17'b01001010001111011,
    17'b01001000101110001,
    17'b01000110001010010,
    17'b01000100011110110,
    17'b01000100111000011,
    17'b01000110001111011,
    17'b01000101100110011,
    17'b01000100000000000,
    17'b01000011010111000,
    17'b01000011000111101,
    17'b01000000011110110,
    17'b00111011110000101,
    17'b00111000011001101,
    17'b00110110011110110,
    17'b00110101000010100,
    17'b00110010111101100,
    17'b00110001010001111,
    17'b00110001110101110,
    17'b00110100001010010,
    17'b00111000100011111,
    17'b00110101111010111,
    17'b00110010111000011,
    17'b00110010100011111,
    17'b00110010011110110,
    17'b00110001100110011,
    17'b00101101000111101,
    17'b00100111100110011,
    17'b00100101010111000,
    17'b00100100100011111,
    17'b00100110111101100,
    17'b00100111001100110,
    17'b00100100100011111,
    17'b00100011000111101,
    17'b00100110011110110,
    17'b00100110100011111,
    17'b00100101000111101,
    17'b00100011100110011,
    17'b00100010111000011,
    17'b00100011011100001,
    17'b00011110000000000,
    17'b00010011101011100,
    17'b00001110000101001,
    17'b00010001010111000,
    17'b00011011001100110,
    17'b00011110111000011,
    17'b00100011101011100,
    17'b00101001000010100,
    17'b00101100010100100,
    17'b00100001010111000,
    17'b00100000001111011,
    17'b00011100000101001,
    17'b00011011100110011,
    17'b00011001000010100,
    17'b00011100011110110,
    17'b00100011010001111,
    17'b00100101000111101,
    17'b00010100011110110,
    17'b00100011000111101,
    17'b00110000111000011,
    17'b00101010101110001,
    17'b00100011011100001,
    17'b00100000010100100,
    17'b00011000110011010,
    17'b00001111010111000,
    17'b00001101100001010,
    17'b00010011010111000,
    17'b00011011100001010,
    17'b00011001000010100,
    17'b00010011001100110,
    17'b00001111110101110,
    17'b00001101110101110,
    17'b00000110000101001,
    17'b00000010010100100,
    17'b00000101111010111,
    17'b00001100011001101,
    17'b00010010001010010,
    17'b00010010101110001,
    17'b00010001100110011,
    17'b00010000111101100,
    17'b00001111110000101,
    17'b00001101110000101,
    17'b00001100001010010,
    17'b00001010110011010,
    17'b00001001010111000,
    17'b00000110111101100,
    17'b00000101110000101,
    17'b00000101000010100,
    17'b00000101010111000,
    17'b00000101111010111,
    17'b00000101101011100,
    17'b00000100110011010,
    17'b00000011111010111,
    17'b00000011000111101,
    17'b00000011100001010,
    17'b00000011010001111,
    17'b00000100001111011,
    17'b00000110011001101,
    17'b00001000110011010,
    17'b00001010100011111,
    17'b00001011001100110,
    17'b00001100000101001,
    17'b00001100010100100,
    17'b00001101000111101,
    17'b00001100100011111,
    17'b00001010110011010,
    17'b00001001010001111,
    17'b00001000011001101,
    17'b00001000001010010,
    17'b00001000011001101,
    17'b00001010010100100,
    17'b00001100000000000,
    17'b00001101110101110,
    17'b00001101000010100,
    17'b00001101100001010,
    17'b00001110111101100,
    17'b00001111100001010,
    17'b00001111110101110,
    17'b00001111110000101,
    17'b00001111101011100,
    17'b00001111000010100,
    17'b00001111000010100,
    17'b00010000011110110,
    17'b00010000110011010,
    17'b00001110010100100,
    17'b00001010000101001,
    17'b00000111011100001,
    17'b00000110010100100,
    17'b00000110001111011,
    17'b00000101100110011,
    17'b00000111000010100,
    17'b00001001110000101,
    17'b00001100011110110,
    17'b00001101111010111,
    17'b00010000100011111,
    17'b00010011100110011,
    17'b00010011100001010,
    17'b00001101101011100,
    17'b00010000110011010,
    17'b00001110110011010,
    17'b00001000111000011,
    17'b00001011001100110,
    17'b00001110100011111,
    17'b00001111000111101,
    17'b00010001110101110,
    17'b00010000100011111,
    17'b00001111110101110,
    17'b00001110001010010,
    17'b00010011000010100,
    17'b00001100111101100,
    17'b00001001100110011,
    17'b11110110110011010,
    17'b11111111100110011,
    17'b00001001010001111,
    17'b11111001100001010,
    17'b11101111001100110,
    17'b11110010101001000,
    17'b11110100011001101,
    17'b11111001010001111,
    17'b11111110110011010,
    17'b00000001001100110,
    17'b00000001010111000,
    17'b11111111111010111,
    17'b00000001100110011,
    17'b00000010010100100,
    17'b00000000001010010,
    17'b11111101110101110,
    17'b11111100011001101,
    17'b11111101000111101,
    17'b11111111100110011,
    17'b00000001100110011,
    17'b00000010011001101,
    17'b00000001011100001,
    17'b11111110110011010,
    17'b11111100100011111,
    17'b11111010110011010,
    17'b11111001111010111,
    17'b11111001101011100,
    17'b11111010010100100,
    17'b11111010100011111,
    17'b11111010001010010,
    17'b11111010011110110,
    17'b11111101011100001,
    17'b00000000100011111,
    17'b00000001110000101,
    17'b00000001111010111,
    17'b00001110111101100,
    17'b00010101001100110,
    17'b00010100000000000,
    17'b00010001110101110,
    17'b00001010110011010,
    17'b00001010100011111,
    17'b00001101101011100,
    17'b00001010000101001,
    17'b00000011000010100,
    17'b00000001101011100,
    17'b11111111111010111,
    17'b00000000011110110,
    17'b00000000000101001,
    17'b00000001000111101,
    17'b11111101110000101,
    17'b00000000100011111,
    17'b00000100100011111,
    17'b00000111100001010,
    17'b00001011111010111,
    17'b00001101110000101,
    17'b00001111000111101,
    17'b00001110111101100,
    17'b00001111000111101,
    17'b00010000000101001,
    17'b00010000101110001,
    17'b00001100001111011,
    17'b00001010110011010,
    17'b00001001000010100,
    17'b00001001100001010,
    17'b00001010111000011,
    17'b00001100001111011,
    17'b00001100101110001,
    17'b00001101100110011,
    17'b00001110010100100,
    17'b00010001011100001,
    17'b00010011100001010,
    17'b00100111101011100,
    17'b00100011100110011,
    17'b00011100101110001,
    17'b00011001001100110,
    17'b00010110111101100,
    17'b00010100111000011,
    17'b00010011001100110,
    17'b00010001001100110,
    17'b00001111100001010,
    17'b00010100011110110,
    17'b00011011010111000,
    17'b00011110101110001,
    17'b00100001000010100,
    17'b00100010000101001,
    17'b00100010001111011,
    17'b00100010011110110,
    17'b00100010001111011,
    17'b00100010101110001,
    17'b00100100001010010,
    17'b00100110101001000,
    17'b00101001100001010,
    17'b00101010000101001,
    17'b00101011010111000,
    17'b00101101111010111,
    17'b00110001100001010,
    17'b00110100110011010,
    17'b00111011010001111,
    17'b00111110111000011,
    17'b00111111000010100,
    17'b00111101111010111,
    17'b00111011011100001,
    17'b00111000010100100,
    17'b00110110100011111,
    17'b00110101001100110,
    17'b00110100001111011,
    17'b00110100001111011,
    17'b00110011110000101,
    17'b00110011100001010,
    17'b00110011110101110,
    17'b00110100010100100,
    17'b00110101000010100,
    17'b00110110001111011,
    17'b00111000011001101,
    17'b00111011110000101,
    17'b00111110001010010,
    17'b01000000011110110,
    17'b01000010111000011,
    17'b01000101001100110,
    17'b01000111101011100,
    17'b01001000111101100,
    17'b01001001100110011,
    17'b01001001000111101,
    17'b01000110111000011,
    17'b01000100011001101,
    17'b01000011101011100,
    17'b01000100011001101,
    17'b01000011101011100,
    17'b01001001111010111,
    17'b00111101010001111,
    17'b01001010110011010,
    17'b01001010100011111,
    17'b01001000000000000,
    17'b01001000101110001,
    17'b01001010000101001,
    17'b01000111100110011,
    17'b01001000011001101,
    17'b01000110011001101,
    17'b01000100010100100,
    17'b01000101000010100,
    17'b01000101001100110,
    17'b01000001100110011,
    17'b01000001100110011,
    17'b00110001101011100,
    17'b00111001000111101,
    17'b01001101000010100,
    17'b01011001000111101,
    17'b01000011000010100,
    17'b11111000000000000,
    17'b11000010110011010,
    17'b11001100111101100,
    17'b11111111011100001,
    17'b00111001100110011,
    17'b01010110001010010,
    17'b01000000011001101,
    17'b00100101101011100,
    17'b00100110101110001,
    17'b00111011100001010,
    17'b01001011110000101,
    17'b01000101100001010,
    17'b00111101100001010,
    17'b00110100110011010,
    17'b00101000010100100,
    17'b00011100011110110,
    17'b00011000101001000,
    17'b00010111111010111,
    17'b00011000011001101,
    17'b00011001000111101,
    17'b00010111110101110,
    17'b00010101110000101,
    17'b00010010101001000,
    17'b00001111110000101,
    17'b00001010111101100,
    17'b00000111000010100,
    17'b00000100001010010,
    17'b00000001010001111,
    17'b11111110010100100,
    17'b11111100111000011,
    17'b11111101100001010,
    17'b11111100111101100,
    17'b11111110001010010,
    17'b11111100000000000,
    17'b11111110000000000,
    17'b11111100011110110,
    17'b11111110000000000,
    17'b11111110001111011,
    17'b00000000101001000,
    17'b00000000111000011,
    17'b00000010111000011,
    17'b00000011100001010,
    17'b00000100100011111,
    17'b00000101110000101,
    17'b00000100001111011,
    17'b00000100111000011,
    17'b00000110001111011,
    17'b00000111101011100,
    17'b00001010101001000,
    17'b00001110001010010,
    17'b00010001000111101,
    17'b00010011100110011,
    17'b00010100101110001,
    17'b00010101110000101,
    17'b00010110100011111,
    17'b00010111000111101,
    17'b00010111001100110,
    17'b00010111010001111,
    17'b00010110111101100,
    17'b00010110011001101,
    17'b00010101111010111,
    17'b00010101011100001,
    17'b00010100100011111,
    17'b00010100000000000,
    17'b00010011101011100,
    17'b00010011001100110,
    17'b00010010110011010,
    17'b00010010101001000,
    17'b00010010100011111,
    17'b00010010010100100,
    17'b00010001111010111,
    17'b00010001010001111,
    17'b00010001010001111,
    17'b00010001100001010,
    17'b00010010011001101,
    17'b00010011110000101,
    17'b00010110010100100,
    17'b00011000110011010,
    17'b00011011010001111,
    17'b00011101010111000,
    17'b00011111101011100,
    17'b00100000110011010,
    17'b00100001110000101,
    17'b00100010010100100,
    17'b00100011000111101,
    17'b00100011110101110,
    17'b00100100110011010,
    17'b00100101111010111,
    17'b00100111000010100,
    17'b00101000110011010,
    17'b00101001111010111,
    17'b00101001111010111,
    17'b00101001010111000,
    17'b00101001010001111,
    17'b00101001010001111,
    17'b00101001010001111,
    17'b00101010000000000,
    17'b00101000001010010,
    17'b00101000010100100,
    17'b00101000111000011,
    17'b00101011011100001,
    17'b00101001110101110,
    17'b00101100000101001,
    17'b00101101110101110,
    17'b00101110010100100,
    17'b00110011000111101,
    17'b00110100100011111,
    17'b00110010001010010,
    17'b00110001000111101,
    17'b00110001110000101,
    17'b00101101111010111,
    17'b00101101000111101,
    17'b00101100011110110,
    17'b00101100011110110,
    17'b00101110001010010,
    17'b00110000011110110,
    17'b00110011100110011,
    17'b00110110010100100,
    17'b00111001001100110,
    17'b00111101000111101,
    17'b00111111100001010,
    17'b01000001011100001,
    17'b01000011000010100,
    17'b01000100101001000,
    17'b01000100111000011,
    17'b01000100110011010,
    17'b01000100101001000,
    17'b01000100011110110,
    17'b01000100001010010,
    17'b01000011110000101,
    17'b01000011001100110,
    17'b01000010000101001,
    17'b01000000111101100,
    17'b00111111110101110,
    17'b00111111010111000,
    17'b00111110111101100,
    17'b00111110111000011,
    17'b00111111001100110,
    17'b00111111110101110,
    17'b01000001000111101,
    17'b01000010101001000,
    17'b01000100000101001,
    17'b01000101010111000,
    17'b01000110111000011,
    17'b01000111101011100,
    17'b01001000010100100,
    17'b01001000100011111,
    17'b01001000111000011,
    17'b01001000111101100,
    17'b01001000110011010,
    17'b01001000010100100,
    17'b01000111100001010,
    17'b01000111010001111,
    17'b01000111011100001,
    17'b01000111110101110,
    17'b01001000100011111,
    17'b01001001010001111,
    17'b01001001100001010,
    17'b01001001010111000,
    17'b01001000111000011,
    17'b01000110100011111,
    17'b01000000001010010,
    17'b00111100001111011,
    17'b00110110101110001,
    17'b00110011100110011,
    17'b00110011000010100,
    17'b00110010111101100,
    17'b00110100000101001,
    17'b00110101010001111,
    17'b00110101101011100,
    17'b00110100111000011,
    17'b00110010101001000,
    17'b00110000001111011,
    17'b00101101010001111,
    17'b00101001010111000,
    17'b00100110011110110,
    17'b00100011000010100,
    17'b00100000000101001,
    17'b00011100000101001,
    17'b00010111001100110,
    17'b00010100001010010,
    17'b00010001010111000,
    17'b00001110101110001,
    17'b00001100011110110,
    17'b00001011010111000,
    17'b00001010111000011,
    17'b00001010000000000,
    17'b00001000000000000,
    17'b00000101110101110,
    17'b00000010111000011,
    17'b11111110101001000,
    17'b11111010101001000,
    17'b11111000011110110,
    17'b11110110000101001,
    17'b11110011110101110,
    17'b11101101101011100,
    17'b11101010111000011,
    17'b11100110111101100,
    17'b11100011000010100,
    17'b11011110111000011,
    17'b11011100100011111,
    17'b11011001010001111,
    17'b11010101010111000,
    17'b11001010001111011,
    17'b11000110001111011,
    17'b11000010101001000,
    17'b11000000001111011,
    17'b11000000000000000,
    17'b10111111011100001,
    17'b10111110101110001,
    17'b10111101111010111,
    17'b10111100001111011,
    17'b10111011001100110,
    17'b10111010101001000,
    17'b10111100000000000,
    17'b10111100011001101,
    17'b10111111100110011,
    17'b11000010010100100,
    17'b11000010110011010,
    17'b11000011110101110,
    17'b11000100100011111,
    17'b11000100111101100,
    17'b11000101000111101,
    17'b11000100001111011,
    17'b11000011011100001,
    17'b11000010001111011,
    17'b11000000111101100,
    17'b10111111110000101,
    17'b10111100111000011,
    17'b10111010011001101,
    17'b10110111110000101,
    17'b10110101100001010,
    17'b10110010111101100,
    17'b10110000001010010,
    17'b10101101000010100,
    17'b10101010001010010,
    17'b10100111100001010,
    17'b10101000001111011,
    17'b10100100010100100,
    17'b10100010100011111,
    17'b10011100001010010,
    17'b10011100111101100,
    17'b10011100011001101,
    17'b10011110010100100,
    17'b10100011001100110,
    17'b10011111010001111,
    17'b10011100111000011,
    17'b10100100100011111,
    17'b10101000100011111,
    17'b10101010011110110,
    17'b10101010111000011,
    17'b10110000100011111,
    17'b10110011110000101,
    17'b10110100111101100,
    17'b10111000001111011,
    17'b10111011111010111,
    17'b10111110001010010,
    17'b10111111101011100,
    17'b11000000101110001,
    17'b11000100001010010,
    17'b11001010011110110,
    17'b11001011010001111,
    17'b11001011110000101,
    17'b11001100101110001,
    17'b11001101011100001,
    17'b11001101100001010,
    17'b11001101110000101,
    17'b11001110101001000,
    17'b11010000000101001,
    17'b11010010000000000,
    17'b11010011101011100,
    17'b11010101100001010,
    17'b11010111000111101,
    17'b11011000110011010,
    17'b11011010000000000,
    17'b11011011000010100,
    17'b11011011111010111,
    17'b11011100101110001,
    17'b11011100101001000,
    17'b11011100110011010,
    17'b11011101100110011,
    17'b11011110101110001,
    17'b11011110011110110,
    17'b11011110000101001,
    17'b11011111011100001,
    17'b11100001100001010,
    17'b11100011101011100,
    17'b11100101001100110,
    17'b11100110001111011,
    17'b11100111000010100,
    17'b11100111101011100,
    17'b11101000001010010,
    17'b11101000010100100,
    17'b11101000100011111,
    17'b11101001000111101,
    17'b11101001110000101,
    17'b11101001111010111,
    17'b11101001110101110,
    17'b11101010011110110,
    17'b11101011000010100,
    17'b11101001111010111,
    17'b11101001000111101,
    17'b11101000000000000,
    17'b11100111001100110,
    17'b11100110011110110,
    17'b11100110000101001,
    17'b11100111111010111,
    17'b11101001010111000,
    17'b11101000011110110,
    17'b11100111010001111,
    17'b11100110101110001,
    17'b11100101100001010,
    17'b11100100010100100,
    17'b11100100100011111,
    17'b11100100110011010,
    17'b11100101101011100,
    17'b11100111000010100,
    17'b11100111010111000,
    17'b11100111011100001,
    17'b11100111101011100,
    17'b11101000000000000,
    17'b11101000101001000,
    17'b11101001001100110,
    17'b11101010000000000,
    17'b11101010010100100,
    17'b11101010101110001,
    17'b11101010101110001,
    17'b11101010111101100,
    17'b11101011001100110,
    17'b11101010101110001,
    17'b11101001110101110,
    17'b11101010000101001,
    17'b11100001010111000,
    17'b11011111000111101,
    17'b11011100011110110,
    17'b11011010001010010,
    17'b11011000000000000,
    17'b11010100100011111,
    17'b11010010101001000,
    17'b11000101110000101,
    17'b10101100100011111,
    17'b10111011000010100,
    17'b11001000011001101,
    17'b11001111000010100,
    17'b11010001000010100,
    17'b11010100101001000,
    17'b11010101001100110,
    17'b11010110111000011,
    17'b11011001010001111,
    17'b11010111010001111,
    17'b11010110111101100,
    17'b11011100101110001,
    17'b11010000111000011,
    17'b11010010010100100,
    17'b11010000101001000,
    17'b11001110111101100,
    17'b11001001110000101,
    17'b11000101111010111,
    17'b11000010111000011,
    17'b10111111010001111,
    17'b10111100011001101,
    17'b10111001100001010,
    17'b10110101110000101,
    17'b10110001000111101,
    17'b10101111100110011,
    17'b10101100000101001,
    17'b10011111110000101,
    17'b10011101101011100,
    17'b10011101000010100,
    17'b10011011110000101,
    17'b10011001010111000,
    17'b10011000111101100,
    17'b10011001110101110,
    17'b10011011110000101,
    17'b10011110100011111,
    17'b10100001010001111,
    17'b10100100001111011,
    17'b10100111010001111,
    17'b10101011100001010,
    17'b10101101110000101,
    17'b10101111110000101,
    17'b10110010000000000,
    17'b10110101000010100,
    17'b10110110111000011,
    17'b10110111111010111,
    17'b10111000001010010,
    17'b10110111110101110,
    17'b10110111011100001,
    17'b10110111010111000,
    17'b10111000000000000,
    17'b10111001000111101,
    17'b10111010001111011,
    17'b10111011101011100,
    17'b10111110000101001,
    17'b11000000000000000,
    17'b11000001100110011,
    17'b11000011000010100,
    17'b11000101000111101,
    17'b11000111011100001,
    17'b11001011000010100,
    17'b11001110111101100,
    17'b11010100101110001,
    17'b11011001001100110,
    17'b11011110010100100,
    17'b11100011001100110,
    17'b11100111110000101,
    17'b11101001000111101,
    17'b11101010101001000,
    17'b11101101010111000,
    17'b11110000100011111,
    17'b11110010100011111,
    17'b11110100001010010,
    17'b11110110001111011,
    17'b11110111111010111,
    17'b11111001011100001,
    17'b11111011010001111,
    17'b11111100001010010,
    17'b11111100101110001,
    17'b11111011101011100,
    17'b11111100011001101,
    17'b11111101011100001,
    17'b11111101100110011,
    17'b11111110110011010,
    17'b00000000101001000,
    17'b00000001101011100,
    17'b00000011100001010,
    17'b00000100000000000,
    17'b00000001110101110,
    17'b00000000111101100,
    17'b00000001100110011,
    17'b00000101001100110,
    17'b00001000011110110,
    17'b00001100001111011,
    17'b00001111110101110,
    17'b00010100101110001,
    17'b00010111111010111,
    17'b00011010101001000,
    17'b00011100111101100,
    17'b00011110101001000,
    17'b00100000100011111,
    17'b00100011000010100,
    17'b00100101000111101,
    17'b00100110111101100,
    17'b00101000100011111,
    17'b00101101000111101,
    17'b00110001010111000,
    17'b00110011110000101,
    17'b00110101000111101,
    17'b00110110100011111,
    17'b00111000010100100,
    17'b00111001000111101,
    17'b00111010110011010,
    17'b00111101111010111,
    17'b01000000001111011,
    17'b01000000101110001,
    17'b01000001001100110,
    17'b01000001111010111,
    17'b01000011000010100,
    17'b01000100000101001,
    17'b01000100001111011,
    17'b01000100001010010,
    17'b01000011100110011,
    17'b01000010100011111,
    17'b01000001100110011,
    17'b01000000100011111,
    17'b00111111100110011,
    17'b00111110001111011,
    17'b00111101010111000,
    17'b00111100011001101,
    17'b00111011011100001,
    17'b00111010110011010,
    17'b00111010011001101,
    17'b00111010000101001,
    17'b00111001101011100,
    17'b00111001000010100,
    17'b00111000101001000,
    17'b00110111011100001,
    17'b00111000001010010,
    17'b00110011010001111,
    17'b00110110110011010,
    17'b00110101101011100,
    17'b00101011100110011,
    17'b00101010001111011,
    17'b00100111000010100,
    17'b00110000011110110,
    17'b00111010101110001,
    17'b01000100000101001,
    17'b01000111000111101,
    17'b01001110001111011,
    17'b01001100111000011,
    17'b01001100011001101,
    17'b01000110101110001,
    17'b01001001110000101,
    17'b01001011110101110,
    17'b01001011110000101,
    17'b01001010110011010,
    17'b01001001100110011,
    17'b01001001010001111,
    17'b01001001110101110,
    17'b01001001100001010,
    17'b01001000011110110,
    17'b01000111010111000,
    17'b01000110001111011,
    17'b01000100000000000,
    17'b01000010010100100,
    17'b01000000000101001,
    17'b00111110111101100,
    17'b00111111010001111,
    17'b00111101000010100,
    17'b00111010110011010,
    17'b00111010101001000,
    17'b00111001011100001,
    17'b00111010110011010,
    17'b00111110000101001,
    17'b01000001110101110,
    17'b01000010111101100,
    17'b00111110001010010,
    17'b00111101110101110,
    17'b00111101100110011,
    17'b00111011010001111,
    17'b00111100000101001,
    17'b00111101011100001,
    17'b00111101010001111,
    17'b00111100000101001,
    17'b00111100011001101,
    17'b00111100101001000,
    17'b00111011101011100,
    17'b00111011100110011,
    17'b00111011100001010,
    17'b00111100000000000,
    17'b00111011011100001,
    17'b00111101011100001,
    17'b00111100011001101,
    17'b00111001000111101,
    17'b00111001111010111,
    17'b00111010011001101,
    17'b00111010010100100,
    17'b00111010011110110,
    17'b00111010011110110,
    17'b00111010011001101,
    17'b00111010011001101,
    17'b00111010101110001,
    17'b00111011010001111,
    17'b00111011111010111,
    17'b00111100011110110,
    17'b00111100101001000,
    17'b00111100111101100,
    17'b00111011101011100,
    17'b00110110101110001,
    17'b00110110101001000,
    17'b00111010111101100,
    17'b00111000101001000,
    17'b00111001110000101,
    17'b00111010011001101,
    17'b01000001011100001,
    17'b01000101010001111,
    17'b01000010001010010,
    17'b01000111100001010,
    17'b01000110011110110,
    17'b01000100111000011,
    17'b01000110101001000,
    17'b01000100001010010,
    17'b01000101100110011,
    17'b01000100110011010,
    17'b01000110101110001,
    17'b01000101010001111,
    17'b01000101100110011,
    17'b01000101011100001,
    17'b01000111110000101,
    17'b01000110011001101,
    17'b01000101010001111,
    17'b01000101101011100,
    17'b01000101000111101,
    17'b01000101000111101,
    17'b01000101011100001,
    17'b01000101000010100,
    17'b01000011011100001,
    17'b01000010100011111,
    17'b01000010101001000,
    17'b01000001011100001,
    17'b01000001001100110,
    17'b01000001100001010,
    17'b01000110111101100,
    17'b01001000101110001,
    17'b01001010010100100,
    17'b01001011110000101,
    17'b01001101010001111,
    17'b01001110000101001,
    17'b01001110000000000,
    17'b01010000000000000,
    17'b01010010001010010,
    17'b01010100001010010,
    17'b01010101010001111,
    17'b01010011100001010,
    17'b01010010011001101,
    17'b01010001111010111,
    17'b01010010111101100,
    17'b01001110101001000,
    17'b01001111000111101,
    17'b01001111110000101,
    17'b01010000100011111,
    17'b01010010111000011,
    17'b01010010001111011,
    17'b01001101000111101,
    17'b01001011000111101,
    17'b01001000111101100,
    17'b01001000010100100,
    17'b01001001000111101,
    17'b01001001110101110,
    17'b01000111011100001,
    17'b01000110011110110,
    17'b01000101100001010,
    17'b01000100111101100,
    17'b01000101000010100,
    17'b01000100111101100,
    17'b01000100101110001,
    17'b01000011100110011,
    17'b01000010100011111,
    17'b01000001010001111,
    17'b01000000001111011,
    17'b00111110110011010,
    17'b00111110001111011,
    17'b00111110000000000,
    17'b00111110101110001,
    17'b00111111101011100,
    17'b00111111101011100,
    17'b00111110111000011,
    17'b00111110001111011,
    17'b00111111011100001,
    17'b01000001011100001,
    17'b01000100000101001,
    17'b01000110101001000,
    17'b01001001000111101,
    17'b01001001100110011,
    17'b01001001011100001,
    17'b01001000101110001,
    17'b01000110111101100,
    17'b01000100001111011,
    17'b01000010101001000,
    17'b01000001001100110,
    17'b01000000000000000,
    17'b00111111010111000,
    17'b00111110110011010,
    17'b00111101101011100,
    17'b00111100010100100,
    17'b00111010000101001,
    17'b00110110000101001,
    17'b00110011100001010,
    17'b00110001110101110,
    17'b00110001000010100,
    17'b00110001000111101,
    17'b00110001000111101,
    17'b00110001000010100,
    17'b00110000110011010,
    17'b00110000000000000,
    17'b00101000000101001,
    17'b00100100111000011,
    17'b00011110101110001,
    17'b00011001100001010,
    17'b00010101010001111,
    17'b00010101000111101,
    17'b00010101110101110,
    17'b00010101111010111,
    17'b00010111110000101,
    17'b00011010000101001,
    17'b00011010111101100,
    17'b00011011010001111,
    17'b00011010101110001,
    17'b00011010010100100,
    17'b00011010000000000,
    17'b00011010000000000,
    17'b00011001110000101,
    17'b00011001110000101,
    17'b00011001110000101,
    17'b00011001100110011,
    17'b00011000100011111,
    17'b00010110111101100,
    17'b00010101010001111,
    17'b00010011010001111,
    17'b00001111110101110,
    17'b00001101010111000,
    17'b00001010111000011,
    17'b00001000011001101,
    17'b00000100110011010,
    17'b00000010000000000,
    17'b11111111110000101,
    17'b11111100111101100,
    17'b11111001100110011,
    17'b11110111110000101,
    17'b11110110001010010,
    17'b11110100010100100,
    17'b11110000011110110,
    17'b11101101100001010,
    17'b11101010011110110,
    17'b11100111100001010,
    17'b11100100001111011,
    17'b11100010001111011,
    17'b11100000100011111,
    17'b11011111000010100,
    17'b11011101011100001,
    17'b11011100011110110,
    17'b11011011110000101,
    17'b11011010111000011,
    17'b11011000111000011,
    17'b11010111100001010,
    17'b11010101011100001,
    17'b11010011001100110,
    17'b11010000011001101,
    17'b11001110111000011,
    17'b11001101001100110,
    17'b11001011100001010,
    17'b11001011010111000,
    17'b11001011000010100,
    17'b11001011001100110,
    17'b11001010111101100,
    17'b11001010001111011,
    17'b11001010000000000,
    17'b11001001011100001,
    17'b11001000010100100,
    17'b11000111011100001,
    17'b11000111001100110,
    17'b11000111011100001,
    17'b11000110111101100,
    17'b11000101010111000,
    17'b11000011011100001,
    17'b11000001100001010,
    17'b10111111011100001,
    17'b10111100101110001,
    17'b10111001111010111,
    17'b10111000011110110,
    17'b10110110101001000,
    17'b10110011110101110,
    17'b10110011000111101,
    17'b10110011000010100,
    17'b10110011000111101,
    17'b10110011011100001,
    17'b10110011101011100,
    17'b10110100001111011,
    17'b10110101001100110,
    17'b10110101100001010,
    17'b10110101100001010,
    17'b10110101110000101,
    17'b10110110000000000,
    17'b10110110001111011,
    17'b10110110101001000,
    17'b10110111001100110,
    17'b10111000000000000,
    17'b10111000011110110,
    17'b10111000011110110,
    17'b10110111101011100,
    17'b10110110000101001,
    17'b10110100111000011,
    17'b10110011111010111,
    17'b10110011010111000,
    17'b10110010110011010,
    17'b10110010011001101,
    17'b10110010011110110,
    17'b10110010100011111,
    17'b10110010110011010,
    17'b10110010110011010,
    17'b10110010111101100,
    17'b10110010011001101,
    17'b10101100101001000,
    17'b10101010011110110,
    17'b10100111010111000,
    17'b10011110110011010,
    17'b10011011011100001,
    17'b10100010010100100,
    17'b10100010111000011,
    17'b10100101101011100,
    17'b10100110011001101,
    17'b10100100001010010,
    17'b10100110111000011,
    17'b11001001100001010,
    17'b11001001000010100,
    17'b11001000011110110,
    17'b11000001111010111,
    17'b10111011100001010,
    17'b10111011010111000,
    17'b10111010010100100,
    17'b10110111100110011,
    17'b10110110011001101,
    17'b10110110111000011,
    17'b10110111111010111,
    17'b10111001101011100,
    17'b10111001101011100,
    17'b10111000111101100,
    17'b10111000000000000,
    17'b10110110111101100,
    17'b10110110100011111,
    17'b10110110001111011,
    17'b10110101111010111,
    17'b10110101010001111,
    17'b10110100100011111,
    17'b10110011110000101,
    17'b10110011100001010,
    17'b10110011000111101,
    17'b10110011000111101,
    17'b10110011001100110,
    17'b10110011101011100,
    17'b10110100111000011,
    17'b10110100111000011,
    17'b10110100001111011,
    17'b10110011110101110,
    17'b10110010101001000,
    17'b10110010000000000,
    17'b10110010000101001,
    17'b10110001110101110,
    17'b10110001100110011,
    17'b10110001110101110,
    17'b10110001111010111,
    17'b10110010001111011,
    17'b10110010001111011,
    17'b10110010001010010,
    17'b10110010001111011,
    17'b10110010010100100,
    17'b10110001110101110,
    17'b10110001101011100,
    17'b10110001010001111,
    17'b10101111100001010,
    17'b10101110111000011,
    17'b10101110011110110,
    17'b10101110011110110,
    17'b10101111010001111,
    17'b10110000011001101,
    17'b10110001010001111,
    17'b10110001000111101,
    17'b10110001000010100,
    17'b10110000110011010,
    17'b10110000100011111,
    17'b10110000010100100,
    17'b10110000001111011,
    17'b10110000101110001,
    17'b10110001001100110,
    17'b10110001011100001,
    17'b10110010010100100,
    17'b10110011100001010,
    17'b10110100101110001,
    17'b10110110010100100,
    17'b10111101110000101,
    17'b11000000011110110,
    17'b11000101110101110,
    17'b11001011000010100,
    17'b11010000011110110,
    17'b11010100110011010,
    17'b11011001000111101,
    17'b11011010100011111,
    17'b11011010001010010,
    17'b11010111011100001,
    17'b11010100100011111,
    17'b11010000111000011,
    17'b11001101000111101,
    17'b11000111100001010,
    17'b11000011010111000,
    17'b10111111000010100,
    17'b10111010011110110,
    17'b10110110011001101,
    17'b10110010001111011,
    17'b10110000010100100,
    17'b10101111100001010,
    17'b10101111110101110,
    17'b10110000101110001,
    17'b10110010000000000,
    17'b10110011100110011,
    17'b10110101010111000,
    17'b10110111010001111,
    17'b10111001110000101,
    17'b10111011110000101,
    17'b10111101110000101,
    17'b11000000101001000,
    17'b11000011001100110,
    17'b11000110111000011,
    17'b11001001001100110,
    17'b11001011111010111,
    17'b11001111100110011,
    17'b11010011100110011,
    17'b11011000101001000,
    17'b11011100000101001,
    17'b11011110000000000,
    17'b11011111000010100,
    17'b11011111111010111,
    17'b11100000110011010,
    17'b11100001001100110,
    17'b11100000100011111,
    17'b11011111110101110,
    17'b11011111001100110,
    17'b11011110101110001,
    17'b11011110000000000,
    17'b11011101000111101,
    17'b11011100000000000,
    17'b11011011101011100,
    17'b11011011000010100,
    17'b11011011000010100,
    17'b11011100000000000,
    17'b11011101000010100,
    17'b11011110100011111,
    17'b11011111111010111,
    17'b11100010001010010,
    17'b11100110000101001,
    17'b11101000111101100,
    17'b11101011110101110,
    17'b11101110110011010,
    17'b11110001010111000,
    17'b11110101000010100,
    17'b11110111110101110,
    17'b11111010001010010,
    17'b11111100010100100,
    17'b11111110001010010,
    17'b11111110111000011,
    17'b11111110111101100,
    17'b11111110011110110,
    17'b11111101111010111,
    17'b11111101010111000,
    17'b11111011100110011,
    17'b11111010011110110,
    17'b11111001101011100,
    17'b11111010110011010,
    17'b11111100000000000,
    17'b11111100001010010,
    17'b11111011110000101,
    17'b11111011101011100,
    17'b11111011000111101,
    17'b11111011000010100,
    17'b11111010110011010,
    17'b11111010011110110,
    17'b11111010001010010,
    17'b11111010000101001,
    17'b11111001110101110,
    17'b11111010001111011,
    17'b11111011010111000,
    17'b11111100110011010,
    17'b11111101110000101,
    17'b11111010111101100,
    17'b11110111011100001,
    17'b11111000001111011,
    17'b11111011110101110,
    17'b11111001010001111,
    17'b11111001010001111,
    17'b11111100001111011,
    17'b11111100101110001,
    17'b11111101001100110,
    17'b11111110001111011,
    17'b11111111110000101,
    17'b00000011011100001,
    17'b00000100010100100,
    17'b00000011111010111,
    17'b00000100011110110,
    17'b00000100111101100,
    17'b00000110000000000,
    17'b00000110101110001,
    17'b00000111010111000,
    17'b00001000011110110,
    17'b00001010001111011,
    17'b00001011001100110,
    17'b00001011100110011,
    17'b00001011100001010,
    17'b00001011010111000,
    17'b00001011010001111,
    17'b00001010100011111,
    17'b00001010011110110,
    17'b00001011100110011,
    17'b00001100110011010,
    17'b00001110101110001,
    17'b00010000000101001,
    17'b00010000000101001,
    17'b00001110001111011,
    17'b00001011010111000,
    17'b00001001100001010,
    17'b00001001010001111,
    17'b00001010101001000,
    17'b00001101011100001,
    17'b00010010100011111,
    17'b00010101100110011,
    17'b00010111011100001,
    17'b00010111110101110,
    17'b00010111000111101,
    17'b00010110111000011,
    17'b00010111010111000,
    17'b00011000001010010,
    17'b00011000111000011,
    17'b00011001000111101,
    17'b00011001100110011,
    17'b00011010100011111,
    17'b00011011100110011,
    17'b00011101000111101,
    17'b00011110100011111,
    17'b00010100010100100,
    17'b11111100110011010,
    17'b11101101110000101,
    17'b00001110111000011,
    17'b00010010011110110,
    17'b00010100001111011,
    17'b00010100010100100,
    17'b00010011010001111,
    17'b00010001110101110,
    17'b00010000011110110,
    17'b00001111000111101,
    17'b00001110110011010,
    17'b00001110101001000,
    17'b00001110110011010,
    17'b00001110110011010,
    17'b00001110011110110,
    17'b00001101110000101,
    17'b00001100101110001,
    17'b00001011010111000,
    17'b00001001000010100,
    17'b00000111010001111,
    17'b00000110000101001,
    17'b00000101011100001,
    17'b00000101101011100,
    17'b00000110111000011,
    17'b00001000111000011,
    17'b00001011011100001,
    17'b00001110001111011,
    17'b00010010001010010,
    17'b00010101001100110,
    17'b00010111110101110,
    17'b00011001110000101,
    17'b00011010010100100,
    17'b00011010011001101,
    17'b00011010110011010,
    17'b00011011010111000,
    17'b00011100010100100,
    17'b00011101001100110,
    17'b00011110011110110,
    17'b00011111111010111,
    17'b00100001101011100,
    17'b00100010101001000,
    17'b00100010111000011,
    17'b00100010100011111,
    17'b00100001100001010,
    17'b00100000100011111,
    17'b00011111001100110,
    17'b00011101111010111,
    17'b00011011111010111,
    17'b00011010001111011,
    17'b00011000001010010,
    17'b00010101110101110,
    17'b00010011010001111,
    17'b00001111111010111,
    17'b00001101100001010,
    17'b00001011001100110,
    17'b00001001010001111,
    17'b00000111010001111,
    17'b00000101111010111,
    17'b00000100101110001,
    17'b00000011110101110,
    17'b00000011000010100,
    17'b00000010101110001,
    17'b00000010011110110,
    17'b00000010010100100,
    17'b00000010011001101,
    17'b00000010111101100,
    17'b00000011100110011,
    17'b00000100100011111,
    17'b00000101100110011,
    17'b00000110111000011,
    17'b00000111100110011,
    17'b00001000000000000,
    17'b00001000001111011,
    17'b00001000001010010,
    17'b00000111110101110,
    17'b00000111000010100,
    17'b00000110000000000,
    17'b00000100100011111,
    17'b00000011010001111,
    17'b00000001100110011,
    17'b11110111111010111,
    17'b11110101100110011,
    17'b11110011111010111,
    17'b11110010011110110,
    17'b11110001011100001,
    17'b11110001000010100,
    17'b11110000110011010,
    17'b11110000011001101,
    17'b11110000001010010,
    17'b11110000001010010,
    17'b11110000100011111,
    17'b11110001010001111,
    17'b11110010011001101,
    17'b11110011000111101,
    17'b11110100000101001,
    17'b11110101000111101,
    17'b11110110111000011,
    17'b11111000011001101,
    17'b11111001100001010,
    17'b11111010001010010,
    17'b11111010101001000,
    17'b11111010100011111,
    17'b11111010101110001,
    17'b11111010101001000,
    17'b11111010001111011,
    17'b11111001010001111,
    17'b11111000000000000,
    17'b11110101110000101,
    17'b11110011110101110,
    17'b11110001101011100,
    17'b11101111100110011,
    17'b11101101100110011,
    17'b11101100100011111,
    17'b11101011010111000,
    17'b11101010001111011,
    17'b11101001100001010,
    17'b11101001110000101,
    17'b11101011101011100,
    17'b11101110011001101,
    17'b11101101111010111,
    17'b11101100010100100,
    17'b11101010111101100,
    17'b11101010010100100,
    17'b11101010101001000,
    17'b11101011000010100,
    17'b11101011010111000,
    17'b11101011000111101,
    17'b11101010101001000,
    17'b11101010011110110,
    17'b11101010111000011,
    17'b11101011110000101,
    17'b11101011011100001,
    17'b11101011000010100,
    17'b11101010011001101,
    17'b11101001101011100,
    17'b11101001010001111,
    17'b11101001000010100,
    17'b11101000100011111,
    17'b11101000000101001,
    17'b11100111011100001,
    17'b11100110111000011,
    17'b11100110000000000,
    17'b11100101010111000,
    17'b11100100111000011,
    17'b11100100000101001,
    17'b11100011100001010,
    17'b11100011001100110,
    17'b11100010111101100,
    17'b11100010111000011,
    17'b11100010101001000,
    17'b11100010101110001,
    17'b11100010100011111,
    17'b11100010111101100,
    17'b11100011011100001,
    17'b11100011110101110,
    17'b11100100011110110,
    17'b11100100010100100,
    17'b11100100000101001,
    17'b11100011111010111,
    17'b11100011110000101,
    17'b11100011010111000,
    17'b11100010110011010,
    17'b11100001111010111,
    17'b11100001100001010,
    17'b11100000101110001,
    17'b11100000001010010,
    17'b11011110111101100,
    17'b11011101111010111,
    17'b11011101000111101,
    17'b11011100000101001,
    17'b11011011110000101,
    17'b11011011100110011,
    17'b11011011100001010,
    17'b11011011110000101,
    17'b11011011110101110,
    17'b11011011101011100,
    17'b11011011000010100,
    17'b11011010101110001,
    17'b11011010101110001,
    17'b11011010110011010,
    17'b11011010100011111,
    17'b11011010000101001,
    17'b11011001010111000,
    17'b11011000101110001,
    17'b11010111111010111,
    17'b11010111101011100,
    17'b11010101000111101,
    17'b11010101011100001,
    17'b11010101111010111,
    17'b11010110110011010,
    17'b11011000000000000,
    17'b11011000111101100,
    17'b11011001110101110,
    17'b11011010100011111,
    17'b11011010111000011,
    17'b11011010111000011,
    17'b11011010101110001,
    17'b11011010101110001,
    17'b11011011000111101,
    17'b11011011011100001,
    17'b11011011100001010,
    17'b11011010111000011,
    17'b11011010001111011,
    17'b11011001001100110,
    17'b11011000001111011,
    17'b11010110101110001,
    17'b11010101101011100,
    17'b11010100110011010,
    17'b11010011100001010,
    17'b11010010101110001,
    17'b11010010000000000,
    17'b11010001110000101,
    17'b11010001101011100,
    17'b11010001110000101,
    17'b11010001011100001,
    17'b11010000101001000,
    17'b11001111110101110,
    17'b11010010101110001,
    17'b11010001111010111,
    17'b11010000110011010,
    17'b11010000001010010,
    17'b11001111111010111,
    17'b11001111111010111,
    17'b11010000001111011,
    17'b11010000111000011,
    17'b11010001100110011,
    17'b11010010101110001,
    17'b11010011000111101,
    17'b11010011010111000,
    17'b11010011010111000,
    17'b11010011000010100,
    17'b11010010111000011,
    17'b11010010111000011,
    17'b11010010101110001,
    17'b11010010100011111,
    17'b11010010101001000,
    17'b11010010011110110,
    17'b11010010111101100,
    17'b11010011010111000,
    17'b11010011110000101,
    17'b11010100001010010,
    17'b11010100011110110,
    17'b11010100111101100,
    17'b11010101010111000,
    17'b11010110100011111,
    17'b11010110101110001,
    17'b11010110000101001,
    17'b11010100110011010,
    17'b11001100000101001,
    17'b11001011000111101,
    17'b11001010010100100,
    17'b11001001010001111,
    17'b11001000011110110,
    17'b11000111100110011,
    17'b11000110111000011,
    17'b11000110011110110,
    17'b11000110001111011,
    17'b11000101110101110,
    17'b11000101001100110,
    17'b11000100111101100,
    17'b11000100111000011,
    17'b11000101010111000,
    17'b11000110100011111,
    17'b11000111100110011,
    17'b11001000010100100,
    17'b11001000110011010,
    17'b11001000111101100,
    17'b11001001000010100,
    17'b11001000110011010,
    17'b11001000011001101,
    17'b11000111111010111,
    17'b11000111000111101,
    17'b11000110010100100,
    17'b11000110000101001,
    17'b11000110000000000,
    17'b11000110000000000,
    17'b11000110000101001,
    17'b11000110011110110,
    17'b11001001001100110,
    17'b11001001101011100,
    17'b11001001001100110,
    17'b11001000000101001,
    17'b11000110000101001,
    17'b11000100101110001,
    17'b11000010110011010,
    17'b11000001000111101,
    17'b10111110101001000,
    17'b10111101001100110,
    17'b10111100010100100,
    17'b10111011110101110,
    17'b10111100001010010,
    17'b10111100101110001,
    17'b10111101001100110,
    17'b10111101001100110,
    17'b10111101000010100,
    17'b10111100011001101,
    17'b10111011010111000,
    17'b10111010000101001,
    17'b10111001001100110,
    17'b10111000110011010,
    17'b10111000010100100,
    17'b10111000000000000,
    17'b10110111111010111,
    17'b10111000000101001,
    17'b10111000000101001,
    17'b10111000100011111,
    17'b10111000110011010,
    17'b10111001100001010,
    17'b10111011001100110,
    17'b10111101001100110,
    17'b11000011000111101,
    17'b11000010100011111,
    17'b11000001101011100,
    17'b11000001000010100,
    17'b11000000001111011,
    17'b10111111111010111,
    17'b10111111110000101,
    17'b10111111100001010,
    17'b10111110111101100,
    17'b10111110110011010,
    17'b10111110011110110,
    17'b10111101110101110,
    17'b10111100101110001,
    17'b10111011111010111,
    17'b10111100001111011,
    17'b10111100111000011,
    17'b10111110001010010,
    17'b10111110011001101,
    17'b10111110101110001,
    17'b10111111111010111,
    17'b11000000011110110,
    17'b11000000111101100,
    17'b11000001010111000,
    17'b11000001111010111,
    17'b11000001010111000,
    17'b11000001010111000,
    17'b11000000110011010,
    17'b10111111111010111,
    17'b10111100011110110,
    17'b10111100111000011,
    17'b10111101100110011,
    17'b10111110111101100,
    17'b11000000011001101,
    17'b11000001010001111,
    17'b11000010001111011,
    17'b11000010101001000,
    17'b11000010011110110,
    17'b11000000111101100,
    17'b10111111111010111,
    17'b10111111001100110,
    17'b10111011000111101,
    17'b10111010101110001,
    17'b10111100011001101,
    17'b10111111000010100,
    17'b11000101110000101,
    17'b11000011000111101,
    17'b11000111000010100,
    17'b11001001010111000,
    17'b11001100001111011,
    17'b11010011000010100,
    17'b11001111110101110,
    17'b11010010001111011,
    17'b11010100001010010,
    17'b11010001100001010,
    17'b11001110001111011,
    17'b11010001000010100,
    17'b11010010011110110,
    17'b11010101110101110,
    17'b11010100101001000,
    17'b11010110010100100,
    17'b11010110101001000,
    17'b11010111010001111,
    17'b11010101100110011,
    17'b11010110001111011,
    17'b11010111011100001,
    17'b11011000111000011,
    17'b11011010111101100,
    17'b11011110011110110,
    17'b11100001000010100,
    17'b11100001101011100,
    17'b11100011010001111,
    17'b11100011001100110,
    17'b11100100110011010,
    17'b11100110100011111,
    17'b11100111010001111,
    17'b11101000000000000,
    17'b11100110101001000,
    17'b11100111100110011,
    17'b11101000111101100,
    17'b11101001110000101,
    17'b11101010000101001,
    17'b11100110111101100,
    17'b11100111110000101,
    17'b11101011000010100,
    17'b11101101110101110,
    17'b11101110110011010,
    17'b11101111010001111,
    17'b11101110111101100,
    17'b11110001011100001,
    17'b11110101011100001,
    17'b11110111101011100,
    17'b11111101000010100,
    17'b11111111110101110,
    17'b00000001000111101,
    17'b11111111000111101,
    17'b11111010010100100,
    17'b11110101000111101,
    17'b11110011010001111,
    17'b11110010111101100,
    17'b11110000001111011,
    17'b11110001100001010,
    17'b11110000011110110,
    17'b11110001010111000,
    17'b11110100011001101,
    17'b11110110100011111,
    17'b11111001110101110,
    17'b11111011110000101,
    17'b11111010000101001,
    17'b11111011010111000,
    17'b11111011110000101,
    17'b11111101010111000,
    17'b11111111101011100,
    17'b11111111110000101,
    17'b11111111000111101,
    17'b11111110001111011,
    17'b11111111100110011,
    17'b00000001110101110,
    17'b00000010101110001,
    17'b00000010011001101,
    17'b00000010001010010,
    17'b00000001110101110,
    17'b00000001111010111,
    17'b00000001100110011,
    17'b00000001000111101,
    17'b00000001000010100,
    17'b00000000011001101,
    17'b11111111101011100,
    17'b11111111110000101,
    17'b00000000000000000,
    17'b00000000011001101,
    17'b00000001000111101,
    17'b00000001110000101,
    17'b00000010000000000,
    17'b00000001111010111,
    17'b00000010001111011,
    17'b00000010011110110,
    17'b00000010000101001,
    17'b00000001001100110,
    17'b11111111110000101,
    17'b11111111010001111,
    17'b11111111100001010,
    17'b11111111100110011,
    17'b00000000001111011,
    17'b00000000101001000,
    17'b00000000111000011,
    17'b00000001000010100,
    17'b00000000101110001,
    17'b00000000101001000,
    17'b00000000110011010,
    17'b00000000110011010,
    17'b00000000011001101,
    17'b11111111110101110,
    17'b11111111101011100,
    17'b00000000000000000,
    17'b00000000011110110,
    17'b00000000111000011,
    17'b00000001001100110,
    17'b00000001111010111,
    17'b00000010011110110,
    17'b00000001111010111,
    17'b00000000000101001,
    17'b00000000000101001,
    17'b11111111000010100,
    17'b11111110101110001,
    17'b11111110001010010,
    17'b11111101110101110,
    17'b11111100101110001,
    17'b11111011100110011,
    17'b11111010010100100,
    17'b11111001101011100,
    17'b11111001110101110,
    17'b11111010100011111,
    17'b11111010111000011,
    17'b11111010101001000,
    17'b11111001100001010,
    17'b11111001000111101,
    17'b11111000011001101,
    17'b11110111100110011,
    17'b11110110001111011,
    17'b11110100111000011,
    17'b11110100000000000,
    17'b11110011010001111,
    17'b11110010100011111,
    17'b11110001100001010,
    17'b11110000111101100,
    17'b11110000100011111,
    17'b11101111101011100,
    17'b11101110111101100,
    17'b11101110010100100,
    17'b11101101011100001,
    17'b11101100101110001,
    17'b11101011111010111,
    17'b11101000110011010,
    17'b11100111011100001,
    17'b11100100101001000,
    17'b11100010010100100,
    17'b11100000001111011,
    17'b11011110101001000,
    17'b11011101010111000,
    17'b11011101101011100,
    17'b11011110101110001,
    17'b11011111111010111,
    17'b11100001100001010,
    17'b11100010000000000,
    17'b11100001100110011,
    17'b11100000100011111,
    17'b11011111010111000,
    17'b11011110111000011,
    17'b11011110111000011,
    17'b11011110110011010,
    17'b11011110001010010,
    17'b11011101001100110,
    17'b11011011100110011,
    17'b11011001101011100,
    17'b11010111000010100,
    17'b11010100111000011,
    17'b11010010110011010,
    17'b11010001000111101,
    17'b11001110111101100,
    17'b11001101100001010,
    17'b11001100001111011,
    17'b11001011000010100,
    17'b11001001110101110,
    17'b11001000110011010,
    17'b11001000000101001,
    17'b11000111100001010,
    17'b11000111001100110,
    17'b11000110011110110,
    17'b11000110000101001,
    17'b11000101101011100,
    17'b11000100011110110,
    17'b11000001010111000,
    17'b11000001111010111,
    17'b11000010011110110,
    17'b11000011000010100,
    17'b11000011010111000,
    17'b11000011100110011,
    17'b11000011110000101,
    17'b11000011110000101,
    17'b11000011100110011,
    17'b11000011011100001,
    17'b11000011010001111,
    17'b11000011001100110,
    17'b11000011000010100,
    17'b11000010101110001,
    17'b11000010011001101,
    17'b11000010001010010,
    17'b11000010010100100,
    17'b11000010101001000,
    17'b11000011001100110,
    17'b11000011001100110,
    17'b11000010111000011,
    17'b11000010100011111,
    17'b11000001110000101,
    17'b11000001001100110,
    17'b11000000101001000,
    17'b11000000010100100,
    17'b10111111101011100,
    17'b10111110111101100,
    17'b10111110000101001,
    17'b10111101000111101,
    17'b10111011101011100,
    17'b10111001111010111,
    17'b10111000001111011,
    17'b10110110110011010,
    17'b10110101100110011,
    17'b10110100101001000,
    17'b10110100000000000,
    17'b10110011001100110,
    17'b10110010011110110,
    17'b10110010000101001,
    17'b10110001101011100,
    17'b10110001001100110,
    17'b10110010000000000,
    17'b10110010010100100,
    17'b10110010101110001,
    17'b10110011000010100,
    17'b10110011110101110,
    17'b10110101000111101,
    17'b10110111011100001,
    17'b10111001010001111,
    17'b10111010111101100,
    17'b10111101001100110,
    17'b11000000101110001,
    17'b11000011110101110,
    17'b11000110110011010,
    17'b11001001111010111,
    17'b11001101100110011,
    17'b11010000000000000,
    17'b11010010000000000,
    17'b11010011011100001,
    17'b11010100101001000,
    17'b11010100110011010,
    17'b11010100011001101,
    17'b11010011111010111,
    17'b11010011010111000,
    17'b11010011001100110,
    17'b11010010101110001,
    17'b11010001111010111,
    17'b11010000111101100,
    17'b11010000010100100,
    17'b11001111100110011,
    17'b11001110111000011,
    17'b11001110000000000,
    17'b11001110001010010,
    17'b11001110011001101,
    17'b11001111010001111,
    17'b11010000001010010,
    17'b11010000110011010,
    17'b11010010000101001,
    17'b11010011101011100,
    17'b11010110000101001,
    17'b11010111110000101,
    17'b11011001010111000,
    17'b11011011000010100,
    17'b11011100011001101,
    17'b11011110001111011,
    17'b11011111011100001,
    17'b11100000011001101,
    17'b11100001010001111,
    17'b11100010101001000,
    17'b11100011110000101,
    17'b11100101000010100,
    17'b11100110011110110,
    17'b11101000111101100,
    17'b11101010110011010,
    17'b11101100101110001,
    17'b11101110101110001,
    17'b11110001110101110,
    17'b11111001101011100,
    17'b11111010111101100,
    17'b11111101000010100,
    17'b11111110111101100,
    17'b00000000110011010,
    17'b00000010001010010,
    17'b00000100101110001,
    17'b00000110101001000,
    17'b00001000001111011,
    17'b00001001010111000,
    17'b00001001110101110,
    17'b00001010001010010,
    17'b00001010010100100,
    17'b00001010010100100,
    17'b00001010011110110,
    17'b00001010101110001,
    17'b00001010111000011,
    17'b00001011100001010,
    17'b00001100101001000,
    17'b00001101100001010,
    17'b00001110000000000,
    17'b00001110110011010,
    17'b00010000001111011,
    17'b00010001100001010,
    17'b00010011000010100,
    17'b00010100010100100,
    17'b00010110000101001,
    17'b00011000010100100,
    17'b00011011110000101,
    17'b00011110011110110,
    17'b00100001011100001,
    17'b00100100011110110,
    17'b00100111000111101,
    17'b00101010001010010,
    17'b00101011110000101,
    17'b00101100111101100,
    17'b00101101011100001,
    17'b00101110010100100,
    17'b00101111000010100,
    17'b00101111101011100,
    17'b00101111110000101,
    17'b00101111010001111,
    17'b00101110010100100,
    17'b00101101011100001,
    17'b00101100110011010,
    17'b00101100110011010,
    17'b00101100001010010,
    17'b00101100100011111,
    17'b00101101011100001,
    17'b00101110110011010,
    17'b00110000111000011,
    17'b00110010111101100,
    17'b00110100110011010,
    17'b00110111000010100,
    17'b00111000100011111,
    17'b00111001000111101,
    17'b00111001111010111,
    17'b00111011011100001,
    17'b00111100110011010,
    17'b00111101011100001,
    17'b00111101001100110,
    17'b00111101010111000,
    17'b00111101110101110,
    17'b00111101110000101,
    17'b00111111010111000,
    17'b01000001100110011,
    17'b01000001100001010,
    17'b01000001011100001,
    17'b01000100001010010,
    17'b01000110001111011,
    17'b01000111000111101,
    17'b01000110100011111,
    17'b01000101100001010,
    17'b01000101111010111,
    17'b01000101101011100,
    17'b01000101100001010,
    17'b01000101100001010,
    17'b01000101010001111,
    17'b01000100011001101,
    17'b01000011010001111,
    17'b01000011100110011,
    17'b01000100101110001,
    17'b01000110000101001,
    17'b01000110100011111,
    17'b01000111000111101,
    17'b01001000011110110,
    17'b01001010000000000,
    17'b01001001011100001,
    17'b01001001000010100,
    17'b01001001111010111,
    17'b01001000111000011,
    17'b01000111001100110,
    17'b01000101100001010,
    17'b01000010111000011,
    17'b01000010000101001,
    17'b01000010011110110,
    17'b01000001011100001,
    17'b01000001001100110,
    17'b01000010000101001,
    17'b01000011001100110,
    17'b01000100101001000,
    17'b01000101011100001,
    17'b01000101100110011,
    17'b01000111110000101,
    17'b01001000000101001,
    17'b01000111100110011,
    17'b01001000011110110,
    17'b01000111100110011,
    17'b01000111010111000,
    17'b01000110010100100,
    17'b01001000000101001,
    17'b01000111011100001,
    17'b01000001110101110,
    17'b00111111110101110,
    17'b01000000111101100,
    17'b01000011100110011,
    17'b01000100111000011,
    17'b01000101010111000,
    17'b01000110000000000,
    17'b01000110001111011,
    17'b01000101100001010,
    17'b01000100101110001,
    17'b01000100101110001,
    17'b01000100011001101,
    17'b01000010000101001,
    17'b01000001010111000,
    17'b01000000011110110,
    17'b01000000101110001,
    17'b01000001010001111,
    17'b01000010000101001,
    17'b01000001110101110,
    17'b01000001111010111,
    17'b01000001001100110,
    17'b00111111100110011,
    17'b00111101000111101,
    17'b00111010110011010,
    17'b00110111101011100,
    17'b00110110011110110,
    17'b00110110001010010,
    17'b00111000001010010,
    17'b00111001000111101,
    17'b00111000111000011,
    17'b00110111101011100,
    17'b00110100111000011,
    17'b00110010011001101,
    17'b00110001001100110,
    17'b00101111100110011,
    17'b00110010000000000,
    17'b00110010110011010,
    17'b00110010001111011,
    17'b00110000101001000,
    17'b00101101110000101,
    17'b00101100000101001,
    17'b00101010100011111,
    17'b00101010000101001,
    17'b00101010101110001,
    17'b00101001111010111,
    17'b00101000101001000,
    17'b00100110111000011,
    17'b00100110001010010,
    17'b00100101011100001,
    17'b00100101000111101,
    17'b00100011111010111,
    17'b00100010010100100,
    17'b00100001001100110,
    17'b00011111111010111,
    17'b00011110110011010,
    17'b00011101101011100,
    17'b00011101001100110,
    17'b00011011101011100,
    17'b00011010011001101,
    17'b00011000011001101,
    17'b00010110000000000,
    17'b00010100111000011,
    17'b00010101101011100,
    17'b00010010011110110,
    17'b00010000000000000,
    17'b00001101011100001,
    17'b00001011001100110,
    17'b00001010011110110,
    17'b00001001001100110,
    17'b00001000011001101,
    17'b00000111001100110,
    17'b00000100111000011,
    17'b00000011010111000,
    17'b00000000011001101,
    17'b11111001111010111,
    17'b11110011101011100,
    17'b11110100011001101,
    17'b11110111111010111,
    17'b11111110000101001,
    17'b00000011110000101,
    17'b00010000010100100,
    17'b00001111111010111,
    17'b00001111110101110,
    17'b00001101101011100,
    17'b00001101000010100,
    17'b00001100001111011,
    17'b00001010010100100,
    17'b00001000001010010,
    17'b00000110111101100,
    17'b00000110110011010,
    17'b00000101100001010,
    17'b00000110011001101,
    17'b00000101110101110,
    17'b00000101011100001,
    17'b00000101010111000,
    17'b00000011111010111,
    17'b00000011101011100,
    17'b00000011100001010,
    17'b00000010101110001,
    17'b00000011010111000,
    17'b00000100101110001,
    17'b00000101000010100,
    17'b00000101001100110,
    17'b00000101110000101,
    17'b00000101110101110,
    17'b00000101001100110,
    17'b00000100001111011,
    17'b00000010011110110,
    17'b00000001110101110,
    17'b00000000100011111,
    17'b11111110011001101,
    17'b11111100100011111,
    17'b11111011111010111,
    17'b11111101110000101,
    17'b11111110000101001,
    17'b11111111000010100,
    17'b00000001110101110,
    17'b00000010100011111,
    17'b00000011000111101,
    17'b00000000101110001,
    17'b00000000011001101,
    17'b00000000001111011,
    17'b11111111100110011,
    17'b11111111010001111,
    17'b00000000011001101,
    17'b00000001001100110,
    17'b00000100010100100,
    17'b00000110101110001,
    17'b00001000000000000,
    17'b00001001100110011,
    17'b00001011110101110,
    17'b00001101100110011,
    17'b00001111010111000,
    17'b00001111000010100,
    17'b00010000010100100,
    17'b00010001101011100,
    17'b00010001101011100,
    17'b00010001100001010,
    17'b00010010010100100,
    17'b00010011110101110,
    17'b00010101000010100,
    17'b00010110001111011,
    17'b00011000001111011,
    17'b00010111011100001,
    17'b00010110110011010,
    17'b00010101010001111,
    17'b00010100001111011,
    17'b00010010011001101,
    17'b00001111100001010,
    17'b00010001110101110,
    17'b00010010011110110,
    17'b00010010001111011,
    17'b00010110111101100,
    17'b00011110010100100,
    17'b00011111000010100,
    17'b00100010100011111,
    17'b00100111100001010,
    17'b00101010001010010,
    17'b00101100100011111,
    17'b00101110000000000,
    17'b00101111000111101,
    17'b00110001001100110,
    17'b00110011010111000,
    17'b00110100111101100,
    17'b00110110001111011,
    17'b00110111100110011,
    17'b00111001100001010,
    17'b00111001000111101,
    17'b00111001000010100,
    17'b00111000101001000,
    17'b00110111110101110,
    17'b00110110101001000,
    17'b00110101011100001,
    17'b00110100101110001,
    17'b00110010100011111,
    17'b00110001110000101,
    17'b00110000111101100,
    17'b00110000100011111,
    17'b00110000101110001,
    17'b00110001100110011,
    17'b00110011100001010,
    17'b00110011010111000,
    17'b00110011011100001,
    17'b00110100011001101,
    17'b00110110000101001,
    17'b00110111110000101,
    17'b00111011101011100,
    17'b00111110001111011,
    17'b01000000101110001,
    17'b01000010000101001,
    17'b01000010001010010,
    17'b01000010001010010,
    17'b01000010101110001,
    17'b01000100010100100,
    17'b01000001100001010,
    17'b01000001010001111,
    17'b00111111110000101,
    17'b00111110000101001,
    17'b00111101000010100,
    17'b00111011101011100,
    17'b00111011010111000,
    17'b00111011000010100,
    17'b00111010101110001,
    17'b00111010000101001,
    17'b00110110100011111,
    17'b00110101110101110,
    17'b00110101110000101,
    17'b00110110100011111,
    17'b00110111001100110,
    17'b00111000000101001,
    17'b00111000110011010,
    17'b00111000111101100,
    17'b00111001001100110,
    17'b00111001011100001,
    17'b00111010000101001,
    17'b00111010110011010,
    17'b00111011110101110,
    17'b00111101000111101,
    17'b00111101101011100,
    17'b00111110000000000,
    17'b00111110001010010,
    17'b00111101111010111,
    17'b00111101010111000,
    17'b00111100111000011,
    17'b00111100000000000,
    17'b00111010011001101,
    17'b00111001000111101,
    17'b00111000001010010,
    17'b00110110101110001,
    17'b00110101101011100,
    17'b00110101000111101,
    17'b00110011110000101,
    17'b00110010101110001,
    17'b00110010011110110,
    17'b00110010100011111,
    17'b00110010001010010,
    17'b00110001100001010,
    17'b00110010101001000,
    17'b00110011000010100,
    17'b00111100000101001,
    17'b00111110011110110,
    17'b00111111110101110,
    17'b01000010100011111,
    17'b01000100001111011,
    17'b01000101010001111,
    17'b01000110000101001,
    17'b01000110011110110,
    17'b01000110100011111,
    17'b01000110000101001,
    17'b01000101110000101,
    17'b01000101110000101,
    17'b01000101001100110,
    17'b01000100111000011,
    17'b01000100110011010,
    17'b01000100011110110,
    17'b01000100001111011,
    17'b01000011110101110,
    17'b01000011011100001,
    17'b01000011001100110,
    17'b01000010111101100,
    17'b01000010101110001,
    17'b01000010000000000,
    17'b01000001100110011,
    17'b01000000110011010,
    17'b01000000001111011,
    17'b00111111010001111,
    17'b00111110110011010,
    17'b00111110011001101,
    17'b00111110010100100,
    17'b00111101111010111,
    17'b00111101101011100,
    17'b00111101110000101,
    17'b00111110000000000,
    17'b00111110100011111,
    17'b00111111010001111,
    17'b00111111101011100,
    17'b00111111111010111,
    17'b00111111010111000,
    17'b00111101110000101,
    17'b00111011100110011,
    17'b00111010101001000,
    17'b00111000011001101,
    17'b00111000001010010,
    17'b00111000001111011,
    17'b00111000000000000,
    17'b00110110100011111,
    17'b00110100101110001,
    17'b00110101100110011,
    17'b00110101000111101,
    17'b00110100001010010,
    17'b00110010001111011,
    17'b00110001011100001,
    17'b00110010011110110,
    17'b00110001001100110,
    17'b00110001111010111,
    17'b00110001100001010,
    17'b00101111100110011,
    17'b00101111000010100,
    17'b00101111100110011,
    17'b00110000000000000,
    17'b00101111101011100,
    17'b00110001000010100,
    17'b00101111011100001,
    17'b00101101101011100,
    17'b00101101010111000,
    17'b00101111000010100,
    17'b00101100111000011,
    17'b00110000000101001,
    17'b00101110011110110,
    17'b00101111111010111,
    17'b00111111000111101,
    17'b01001100000000000,
    17'b00111100100011111,
    17'b00111011100001010,
    17'b00101001100001010,
    17'b00011100101001000,
    17'b00010101111010111,
    17'b00010101000010100,
    17'b00100001001100110,
    17'b00100100000000000,
    17'b00100011110000101,
    17'b00100100010100100,
    17'b00100100001111011,
    17'b00100011110000101,
    17'b00100000100011111,
    17'b00100000110011010,
    17'b00011111110000101,
    17'b00100000100011111,
    17'b00011111100001010,
    17'b00011110101110001,
    17'b00011101101011100,
    17'b00011101100110011,
    17'b00011101000111101,
    17'b00011101001100110,
    17'b00011100111101100,
    17'b00011100011110110,
    17'b00011011101011100,
    17'b00011100001010010,
    17'b00011100001111011,
    17'b00011011110101110,
    17'b00011010101001000,
    17'b00011011010001111,
    17'b00011010000000000,
    17'b00011001011100001,
    17'b00011000001111011,
    17'b00011001101011100,
    17'b00011000101110001,
    17'b00010111001100110,
    17'b00011011100110011,
    17'b00011000111000011,
    17'b00010010110011010,
    17'b00010011011100001,
    17'b00001100111101100,
    17'b11111000111000011,
    17'b00001011010001111,
    17'b00001000011001101,
    17'b00000110101001000,
    17'b00000110010100100,
    17'b00000110101110001,
    17'b00000110111101100,
    17'b00000101100001010,
    17'b00000101000010100,
    17'b00000010100011111,
    17'b00000100001111011,
    17'b00000001001100110,
    17'b11111100101001000,
    17'b11111011000010100,
    17'b11111001001100110,
    17'b11111000101110001,
    17'b11111000000000000,
    17'b11111000111101100,
    17'b11111010100011111,
    17'b11111001110101110,
    17'b11111000111101100,
    17'b11110111010111000,
    17'b11110110011001101,
    17'b11110101110101110,
    17'b11111100000000000,
    17'b11111010001010010,
    17'b11111000110011010,
    17'b00010001000111101,
    17'b11111010100011111,
    17'b11101010111000011,
    17'b11101000101110001,
    17'b11101010001010010,
    17'b11101101010001111,
    17'b11110001000010100,
    17'b11110110101001000,
    17'b11110101110000101,
    17'b11110100111000011,
    17'b11110110001111011,
    17'b11111111110101110,
    17'b11111000000101001,
    17'b11110010111000011,
    17'b11110011010001111,
    17'b11111010001010010,
    17'b11111101000111101,
    17'b11110100110011010,
    17'b11110101010111000,
    17'b11111110001111011,
    17'b11110110000000000,
    17'b11111101001100110,
    17'b11110100011001101,
    17'b11110100111101100,
    17'b11111110011001101,
    17'b00000011010001111,
    17'b11110001100001010,
    17'b11101100001111011,
    17'b11101011000010100,
    17'b11101101101011100,
    17'b11101100100011111,
    17'b11101101011100001,
    17'b11101110000000000,
    17'b11101111010001111,
    17'b11101110100011111,
    17'b11101110100011111,
    17'b11101001101011100,
    17'b11100010101110001,
    17'b11100001001100110,
    17'b11011001100110011,
    17'b11010100011001101,
    17'b11010100010100100,
    17'b11010110101001000,
    17'b11011001001100110,
    17'b11010001101011100,
    17'b11001110101110001,
    17'b11001011100001010,
    17'b11001010000101001,
    17'b11001001100001010,
    17'b11001001001100110,
    17'b11000111110101110,
    17'b11001000111101100,
    17'b11001001000111101,
    17'b11001010011110110,
    17'b11001011010001111,
    17'b11001100000101001,
    17'b11001010111000011,
    17'b11001000001111011,
    17'b11000101111010111,
    17'b11000011110000101,
    17'b11000010001010010,
    17'b10111111110101110,
    17'b10111110011001101,
    17'b10111100111000011,
    17'b10111011100001010,
    17'b10111010110011010,
    17'b10111010111101100,
    17'b10111011010111000,
    17'b10111100001010010,
    17'b10111100101110001,
    17'b10111101010111000,
    17'b10111110000000000,
    17'b10111110110011010,
    17'b10111111010001111,
    17'b10111111100001010,
    17'b10111111110000101,
    17'b10111110110011010,
    17'b10111110111000011,
    17'b10111111000111101,
    17'b10111110111000011,
    17'b10111110010100100,
    17'b10111101110000101,
    17'b10111101010001111,
    17'b10111101001100110,
    17'b10111100101110001,
    17'b10111100011110110,
    17'b10111100001010010,
    17'b10111011100110011,
    17'b10111010110011010,
    17'b10111001110000101,
    17'b10111001100110011,
    17'b10111001111010111,
    17'b10111010000101001,
    17'b10111001101011100,
    17'b10111001100110011,
    17'b10111010000000000,
    17'b10111010111101100,
    17'b10111100011110110,
    17'b10111110100011111,
    17'b10111111110000101,
    17'b11000001100001010,
    17'b11000001001100110,
    17'b11000100001010010,
    17'b11000100101110001,
    17'b11000100100011111,
    17'b11000110000101001,
    17'b11000111000010100,
    17'b11000101001100110,
    17'b11000100001111011,
    17'b11000011010001111,
    17'b11000010010100100,
    17'b11000001000111101,
    17'b11000000101001000,
    17'b11000000010100100,
    17'b11000000110011010,
    17'b10111111101011100,
    17'b10111111110000101,
    17'b11000001001100110,
    17'b11000001100001010,
    17'b11000011111010111,
    17'b11000100011110110,
    17'b11000100111000011,
    17'b11000101111010111,
    17'b11001000001010010,
    17'b11001010101110001,
    17'b11001001100110011,
    17'b11001010000000000,
    17'b11001011000010100,
    17'b11001011000111101,
    17'b11000111101011100,
    17'b11001011010111000,
    17'b11001100110011010,
    17'b11010000011001101,
    17'b11010100000101001,
    17'b11010111011100001,
    17'b11011001000010100,
    17'b11011011101011100,
    17'b11011100000000000,
    17'b11011101100110011,
    17'b11011110101110001,
    17'b11100000101001000,
    17'b11100001101011100,
    17'b11100010010100100,
    17'b11100100101001000,
    17'b11100101100110011,
    17'b11100110111000011,
    17'b11100111010001111,
    17'b11100111110101110,
    17'b11101000110011010,
    17'b11101001111010111,
    17'b11101000111101100,
    17'b11101000011001101,
    17'b11101001000111101,
    17'b11101010011110110,
    17'b11101011000111101,
    17'b11101011001100110,
    17'b11101011110000101,
    17'b11101101110000101,
    17'b11101111010111000,
    17'b11110001000010100,
    17'b11110010000101001,
    17'b11110010111000011,
    17'b11110111100110011,
    17'b11111000100011111,
    17'b11111001010111000,
    17'b11111010001111011,
    17'b11111011010001111,
    17'b11111100000101001,
    17'b11111100111101100,
    17'b11111101110000101,
    17'b11111110101001000,
    17'b11111110111101100,
    17'b11111110110011010,
    17'b11111110111000011,
    17'b11111111000111101,
    17'b00000000000101001,
    17'b00000001010001111,
    17'b00000001001100110,
    17'b00000000111000011,
    17'b00000000011001101,
    17'b00000000111000011,
    17'b00000010001010010,
    17'b00000011100110011,
    17'b00000100000101001,
    17'b00000100101110001,
    17'b00000110100011111,
    17'b00001000101110001,
    17'b00001010111101100,
    17'b00001011011100001,
    17'b00001101000010100,
    17'b00001110001111011,
    17'b00001111011100001,
    17'b00001111111010111,
    17'b00010000010100100,
    17'b00010000110011010,
    17'b00010000111000011,
    17'b00010000101110001,
    17'b00010000101110001,
    17'b00010001010111000,
    17'b00010010001010010,
    17'b00010010111000011,
    17'b00010011000010100,
    17'b00010011000010100,
    17'b00010011000010100,
    17'b00010000101110001,
    17'b00001011101011100,
    17'b00001100111000011,
    17'b00001100101110001,
    17'b00001011010111000,
    17'b00001110000101001,
    17'b00010000001010010,
    17'b00010100100011111,
    17'b00010111100001010,
    17'b00011000111000011,
    17'b00011000101110001,
    17'b00010111000111101,
    17'b00010100110011010,
    17'b00010010111101100,
    17'b00010010111000011,
    17'b00001111110101110,
    17'b00010000000000000,
    17'b00001111101011100,
    17'b00001110000000000,
    17'b00001010111101100,
    17'b00001011000010100,
    17'b00001011011100001,
    17'b00001010011110110,
    17'b00000111000010100,
    17'b00000101110000101,
    17'b00000101001100110,
    17'b00000101100001010,
    17'b00000101101011100,
    17'b00000100101001000,
    17'b00000100010100100,
    17'b00000100000101001,
    17'b00000011110101110,
    17'b00000011101011100,
    17'b00000010101110001,
    17'b00000010001010010,
    17'b00000010001111011,
    17'b00000010001111011,
    17'b00000010001010010,
    17'b00000010011110110,
    17'b00000010101110001,
    17'b00000010111000011,
    17'b00000010100011111,
    17'b00000010011110110,
    17'b00000010001010010,
    17'b00000001010111000,
    17'b11111111110000101,
    17'b11110000111000011,
    17'b11101101000010100,
    17'b11101010111000011,
    17'b11101011000111101,
    17'b11110000010100100,
    17'b11110011100110011,
    17'b11111000001010010,
    17'b11111011100110011,
    17'b11111110111101100,
    17'b00000000011001101,
    17'b00000000101110001,
    17'b00000000100011111,
    17'b00000000001111011,
    17'b11111111101011100,
    17'b11111111000010100,
    17'b11111110010100100,
    17'b11111110000101001,
    17'b11111101101011100,
    17'b11111101010111000,
    17'b11111101000111101,
    17'b11111100111000011,
    17'b11111100110011010,
    17'b11111101010111000,
    17'b11111110011110110,
    17'b11111110101001000,
    17'b11111110011110110,
    17'b11111110001010010,
    17'b11111101110000101,
    17'b11111101100110011,
    17'b11111101010001111,
    17'b11111100111000011,
    17'b11111100110011010,
    17'b11111111001100110,
    17'b11111100001010010,
    17'b11111011000111101,
    17'b11111001110000101,
    17'b11111000011110110,
    17'b11110111101011100,
    17'b11110110001010010,
    17'b11110100000101001,
    17'b11110011101011100,
    17'b11110001010001111,
    17'b11110000001111011,
    17'b11101110111000011,
    17'b11101100000000000,
    17'b11101010001111011,
    17'b11101001010001111,
    17'b11100111100001010,
    17'b11101000011001101,
    17'b11101001100001010,
    17'b11101100110011010,
    17'b11101101111010111,
    17'b11101100111101100,
    17'b11101011100110011,
    17'b11101100101110001,
    17'b11101111010111000,
    17'b11110010010100100,
    17'b11111101001100110,
    17'b00000000110011010,
    17'b11111010111101100,
    17'b11110111100001010,
    17'b11111000001010010,
    17'b11110100110011010,
    17'b11110000011001101,
    17'b11101111101011100,
    17'b11110000100011111,
    17'b11101000001010010,
    17'b11101000011001101,
    17'b11101000011110110,
    17'b11101010001111011,
    17'b11100111111010111,
    17'b11100110101110001,
    17'b11100101110000101,
    17'b11100011010001111,
    17'b11100000001111011,
    17'b11011110111101100,
    17'b11011100011001101,
    17'b11011001100110011,
    17'b11010111111010111,
    17'b11011000001010010,
    17'b11010111101011100,
    17'b11010110011001101,
    17'b11010101100110011,
    17'b11010101000010100,
    17'b11010101010111000,
    17'b11010111011100001,
    17'b11011001100110011,
    17'b11011011110101110,
    17'b11011100010100100,
    17'b11011010000000000,
    17'b11011000100011111,
    17'b11011000011110110,
    17'b11011001001100110,
    17'b11011001100001010,
    17'b11011000110011010,
    17'b11010111110000101,
    17'b11010110000101001,
    17'b11010101000010100,
    17'b11010011110000101,
    17'b11010010011110110,
    17'b11010000010100100,
    17'b11001110101110001,
    17'b11001101010111000,
    17'b11001101000010100,
    17'b11001110001010010,
    17'b11001111010001111,
    17'b11001111111010111,
    17'b11010000011110110,
    17'b11010001000010100,
    17'b11010001111010111,
    17'b11010010101001000,
    17'b11010001010111000,
    17'b11001111111010111,
    17'b11001110000101001,
    17'b11001101001100110,
    17'b11001101000111101,
    17'b11001100111101100,
    17'b11001101000010100,
    17'b11001101001100110,
    17'b11001011010111000,
    17'b11001001010111000,
    17'b11000111000010100,
    17'b11001000010100100,
    17'b11001001010001111,
    17'b11001011011100001,
    17'b11001101100110011,
    17'b11010001000010100,
    17'b11010001110101110,
    17'b11010010101001000,
    17'b11010011010001111,
    17'b11010010010100100,
    17'b11010000101110001,
    17'b11001111111010111,
    17'b11001111000010100,
    17'b11001110000101001,
    17'b11001100101110001,
    17'b11001010111101100,
    17'b11001001101011100,
    17'b11001001010001111,
    17'b11001010011110110,
    17'b11001011100110011,
    17'b11001100011110110,
    17'b11001110010100100,
    17'b11001111100110011,
    17'b11010000101001000,
    17'b11010000101110001,
    17'b11001111110101110,
    17'b11001100001111011,
    17'b11001011100001010,
    17'b11001011100001010,
    17'b11001100001010010,
    17'b11001100111101100,
    17'b11001101101011100,
    17'b11001110100011111,
    17'b11001110111000011,
    17'b11001110111000011,
    17'b11001111000111101,
    17'b11001111000010100,
    17'b11001111011100001,
    17'b11001111100110011,
    17'b11010000011001101,
    17'b11010001011100001,
    17'b11010010011110110,
    17'b11010011100110011,
    17'b11010110001111011,
    17'b11010110101110001,
    17'b11010110011001101,
    17'b11010111100110011,
    17'b11011000100011111,
    17'b11011001100001010,
    17'b11011011001100110,
    17'b11011101011100001,
    17'b11011111011100001,
    17'b11100001001100110,
    17'b11100010000000000,
    17'b11100011100001010,
    17'b11100011001100110,
    17'b11100010101001000,
    17'b11100011100001010,
    17'b11100100101001000,
    17'b11100101000010100,
    17'b11100101110000101,
    17'b11100110101001000,
    17'b11101000000000000,
    17'b11101010001010010,
    17'b11101100000000000,
    17'b11101101111010111,
    17'b11101111110101110,
    17'b11110010010100100,
    17'b11110100010100100,
    17'b11110110001010010,
    17'b11111000001111011,
    17'b11111011000010100,
    17'b11111100111101100,
    17'b11111110111101100,
    17'b00000000101110001,
    17'b00000010110011010,
    17'b00000011100110011,
    17'b00000100101001000,
    17'b00000101110000101,
    17'b00000110110011010,
    17'b00000111100001010,
    17'b00001000001010010,
    17'b00001000110011010,
    17'b00001001011100001,
    17'b00001011010111000,
    17'b00001101000111101,
    17'b00001111000111101,
    17'b00010001000010100,
    17'b00010010101110001,
    17'b00010100001111011,
    17'b00010100111000011,
    17'b00010101000111101,
    17'b00010101001100110,
    17'b00010101110101110,
    17'b00010110111101100,
    17'b00011000011001101,
    17'b00011001110000101,
    17'b00011011011100001,
    17'b00011100011001101,
    17'b00011101010001111,
    17'b00011110010100100,
    17'b00011111110000101,
    17'b00100001110000101,
    17'b00100011000111101,
    17'b00100100010100100,
    17'b00100101010111000,
    17'b00100110100011111,
    17'b00100111010111000,
    17'b00101000101110001
};

parameter logic signed [`ACC_WIDTH-1:0] AZ_TEST_VECTOR[`NUM_ELEMENTS] = {
    17'b00011000011110110,
    17'b00011000110011010,
    17'b00011001010001111,
    17'b00011001111010111,
    17'b00011010011110110,
    17'b00011011000111101,
    17'b00011011101011100,
    17'b00011100101001000,
    17'b00011101100001010,
    17'b00011110011110110,
    17'b00011111001100110,
    17'b00011111010111000,
    17'b00011111100110011,
    17'b00011111110000101,
    17'b00011111110000101,
    17'b00011111110000101,
    17'b00011111101011100,
    17'b00100000000000000,
    17'b00100000011001101,
    17'b00100001010001111,
    17'b00100001111010111,
    17'b00100011010001111,
    17'b00100100100011111,
    17'b00100110010100100,
    17'b00101000000101001,
    17'b00101010100011111,
    17'b00101100100011111,
    17'b00101110100011111,
    17'b00110000001111011,
    17'b00110010001111011,
    17'b00110011010001111,
    17'b00110100001111011,
    17'b00110100111101100,
    17'b00110100110011010,
    17'b00110100100011111,
    17'b00110100011001101,
    17'b00110011000111101,
    17'b00110010110011010,
    17'b00110011100001010,
    17'b00110100111101100,
    17'b00110111100001010,
    17'b00111001000111101,
    17'b00111001101011100,
    17'b00111001000111101,
    17'b00110111000111101,
    17'b00110101100001010,
    17'b00110100001010010,
    17'b00110011010001111,
    17'b00110010010100100,
    17'b00110001111010111,
    17'b00110001101011100,
    17'b00110001010111000,
    17'b00110001001100110,
    17'b00110000110011010,
    17'b00110000101001000,
    17'b00110000101001000,
    17'b00110000110011010,
    17'b00110001010001111,
    17'b00110001101011100,
    17'b00110010101110001,
    17'b00110100000000000,
    17'b00110101011100001,
    17'b00110110110011010,
    17'b00111000100011111,
    17'b00111000100011111,
    17'b00110101111010111,
    17'b00110010110011010,
    17'b00101110110011010,
    17'b00101011101011100,
    17'b00101001001100110,
    17'b00101000111000011,
    17'b00101010101110001,
    17'b00101101110101110,
    17'b00110001110000101,
    17'b00110100111000011,
    17'b00110011100110011,
    17'b00101000011001101,
    17'b00100001110000101,
    17'b00010110001111011,
    17'b00001010111101100,
    17'b00000100011110110,
    17'b00010000000000000,
    17'b00100001000111101,
    17'b00111010101001000,
    17'b01010110010100100,
    17'b01101110111101100,
    17'b01110011110000101,
    17'b01101101110000101,
    17'b01011111001100110,
    17'b01000111010111000,
    17'b00110101011100001,
    17'b00100111000010100,
    17'b00011101101011100,
    17'b00011001000010100,
    17'b00011001111010111,
    17'b00011101100110011,
    17'b00100010000101001,
    17'b00100110111101100,
    17'b00101001000010100,
    17'b00101010000000000,
    17'b00101011100001010,
    17'b00101011011100001,
    17'b00101010010100100,
    17'b00101000100011111,
    17'b00101000100011111,
    17'b00101001010111000,
    17'b00101011001100110,
    17'b00101110001010010,
    17'b00110000000000000,
    17'b00110000110011010,
    17'b00110001110000101,
    17'b00110000011001101,
    17'b00101101110101110,
    17'b00101011010111000,
    17'b00101001011100001,
    17'b00101000011001101,
    17'b00101000101110001,
    17'b00101010000000000,
    17'b00101011111010111,
    17'b00101110111000011,
    17'b00110001001100110,
    17'b00110101011100001,
    17'b00111010101110001,
    17'b00111000001010010,
    17'b00110010000000000,
    17'b00110001010111000,
    17'b00110001110101110,
    17'b00110000101001000,
    17'b00101101010001111,
    17'b00101100001111011,
    17'b00101011000010100,
    17'b00101010001010010,
    17'b00101001000010100,
    17'b00101000111000011,
    17'b00101001010111000,
    17'b00101001000010100,
    17'b00101000000101001,
    17'b00100110000000000,
    17'b00100100011001101,
    17'b00100001000010100,
    17'b00011110111101100,
    17'b00011111001100110,
    17'b00100001000111101,
    17'b00100010011001101,
    17'b00100011100110011,
    17'b00100010011001101,
    17'b00100011011100001,
    17'b00100101001100110,
    17'b00100111100001010,
    17'b00101010000101001,
    17'b00101010101001000,
    17'b00101001000010100,
    17'b00101000010100100,
    17'b00100111111010111,
    17'b00100110011110110,
    17'b00100111010111000,
    17'b00100111010001111,
    17'b00101001001100110,
    17'b00101010001111011,
    17'b00101011000111101,
    17'b00101011010001111,
    17'b00101011010001111,
    17'b00101011011100001,
    17'b00101011111010111,
    17'b00101100010100100,
    17'b00101011100110011,
    17'b00101011110101110,
    17'b00101010111000011,
    17'b00101000110011010,
    17'b00101000001111011,
    17'b00101000101001000,
    17'b00101000100011111,
    17'b00101000000000000,
    17'b00101000010100100,
    17'b00101000111000011,
    17'b00101010010100100,
    17'b00110010101110001,
    17'b00110000001010010,
    17'b00101110000101001,
    17'b00101100111000011,
    17'b00101001010111000,
    17'b00100111111010111,
    17'b00100001110101110,
    17'b00100100000101001,
    17'b00100100011001101,
    17'b00011010100011111,
    17'b00001111001100110,
    17'b00000000011110110,
    17'b11101100111101100,
    17'b11101100000101001,
    17'b11110011101011100,
    17'b11111111100110011,
    17'b00001110111000011,
    17'b00011000101110001,
    17'b00100000001111011,
    17'b00100101010111000,
    17'b00101001000111101,
    17'b00101011100001010,
    17'b00101110110011010,
    17'b00110010011110110,
    17'b00111010011001101,
    17'b00111100111000011,
    17'b00110111010111000,
    17'b00110100110011010,
    17'b00110100010100100,
    17'b00101011010111000,
    17'b00100001101011100,
    17'b00011101111010111,
    17'b00010111010001111,
    17'b00010011010001111,
    17'b00010001100110011,
    17'b00010010011001101,
    17'b00010100111101100,
    17'b00011010111101100,
    17'b00100001010001111,
    17'b00101000101001000,
    17'b00110000000101001,
    17'b00111011000010100,
    17'b01000011110000101,
    17'b01001100000101001,
    17'b01010011011100001,
    17'b01011010111000011,
    17'b01011101111010111,
    17'b01011110100011111,
    17'b01011100100011111,
    17'b01010111110000101,
    17'b01001110011110110,
    17'b01000110101001000,
    17'b00111110111000011,
    17'b00110111110000101,
    17'b00101111110101110,
    17'b00101011011100001,
    17'b00100111110101110,
    17'b00100100111000011,
    17'b00100001100110011,
    17'b00011111100001010,
    17'b00011101111010111,
    17'b00011100001111011,
    17'b00011011011100001,
    17'b00011011000111101,
    17'b00011011000010100,
    17'b00011011001100110,
    17'b00011100000101001,
    17'b00011101101011100,
    17'b00011110011001101,
    17'b00010100100011111,
    17'b00001101110101110,
    17'b00100101110000101,
    17'b01001101111010111,
    17'b00101010000000000,
    17'b00010110111000011,
    17'b00011111011100001,
    17'b00101111011100001,
    17'b00100110011110110,
    17'b01000110011001101,
    17'b00110000011001101,
    17'b00100111001100110,
    17'b00100110101110001,
    17'b00101001101011100,
    17'b00100100011001101,
    17'b00100101100110011,
    17'b00100011110101110,
    17'b00100100111101100,
    17'b00100011110000101,
    17'b00100010111000011,
    17'b00100101100001010,
    17'b00100110101110001,
    17'b00100101011100001,
    17'b00100101100001010,
    17'b00100110011001101,
    17'b00100100011001101,
    17'b00100111010111000,
    17'b00100110110011010,
    17'b00100110011110110,
    17'b00100110110011010,
    17'b00100110101001000,
    17'b00100111110000101,
    17'b00100101000111101,
    17'b00100101100110011,
    17'b00100101111010111,
    17'b00100111000111101,
    17'b00100111110101110,
    17'b00100101111010111,
    17'b00100010111101100,
    17'b00100011111010111,
    17'b00100100001111011,
    17'b00100110111000011,
    17'b00100110100011111,
    17'b00100110100011111,
    17'b00100110011110110,
    17'b00100110011001101,
    17'b00100110000000000,
    17'b00100110000000000,
    17'b00100110010100100,
    17'b00100110001010010,
    17'b00100110001010010,
    17'b00100110001010010,
    17'b00100110001010010,
    17'b00100110000101001,
    17'b00100110001010010,
    17'b00100110000000000,
    17'b00100110000101001,
    17'b00100110000000000,
    17'b00100110000000000,
    17'b00100110000000000,
    17'b00100110000000000,
    17'b00100101110101110,
    17'b00100101110101110,
    17'b00100101111010111,
    17'b00100101111010111,
    17'b00100110000000000,
    17'b00100110000000000,
    17'b00100101110101110,
    17'b00100101111010111,
    17'b00100110000101001,
    17'b00100110000101001,
    17'b00100110001111011,
    17'b00100110001111011,
    17'b00100110011001101,
    17'b00100110010100100,
    17'b00100110001111011,
    17'b00100110001010010,
    17'b00100110001111011,
    17'b00100110001010010,
    17'b00100110001010010,
    17'b00100110001010010,
    17'b00100110000101001,
    17'b00100110000101001,
    17'b00100110000101001,
    17'b00100110000101001,
    17'b00100110000101001,
    17'b00100110000101001,
    17'b00100110001010010,
    17'b00100110001010010,
    17'b00100110001111011,
    17'b00100110001111011,
    17'b00100110000000000,
    17'b00100110001010010,
    17'b00100110001010010,
    17'b00100110001111011,
    17'b00100110010100100,
    17'b00100110011110110,
    17'b00100110011110110,
    17'b00100110001111011,
    17'b00100110011001101,
    17'b00100110100011111,
    17'b00100110011001101,
    17'b00100110001010010,
    17'b00100110000101001,
    17'b00100110001010010,
    17'b00100110001111011,
    17'b00100110010100100,
    17'b00100110011001101,
    17'b00100110011110110,
    17'b00100110011001101,
    17'b00100110001010010,
    17'b00100110000101001,
    17'b00100110001111011,
    17'b00100110001111011,
    17'b00100110001111011,
    17'b00100110001111011,
    17'b00100110001010010,
    17'b00100110001010010,
    17'b00100110001111011,
    17'b00100101111010111,
    17'b00100100000000000,
    17'b00100001010111000,
    17'b00100010100011111,
    17'b00100101100001010,
    17'b00100111011100001,
    17'b00101000111101100,
    17'b00101010001111011,
    17'b00101001000010100,
    17'b00100110011001101,
    17'b00101000100011111,
    17'b00100101011100001,
    17'b00100101101011100,
    17'b00100110001010010,
    17'b00100111001100110,
    17'b00100110101110001,
    17'b00100101110000101,
    17'b00100101001100110,
    17'b00100100101110001,
    17'b00100110001111011,
    17'b00100110101110001,
    17'b00100111001100110,
    17'b00100111011100001,
    17'b00100110111101100,
    17'b00100101110000101,
    17'b00100101111010111,
    17'b00100101111010111,
    17'b00100101110101110,
    17'b00100110111000011,
    17'b00100110100011111,
    17'b00100110000000000,
    17'b00100101100001010,
    17'b00100101100001010,
    17'b00100101110101110,
    17'b00100110011110110,
    17'b00100110110011010,
    17'b00100110111000011,
    17'b00100110111000011,
    17'b00100110111101100,
    17'b00100110110011010,
    17'b00100110110011010,
    17'b00101000110011010,
    17'b00110000111101100,
    17'b00111100111000011,
    17'b00110011110101110,
    17'b00100101100001010,
    17'b00100100101110001,
    17'b00011110111000011,
    17'b00101010001111011,
    17'b00111000101001000,
    17'b00110011001100110,
    17'b00101110001010010,
    17'b00101101110101110,
    17'b00100110111101100,
    17'b00101101001100110,
    17'b00101100111101100,
    17'b00100010101001000,
    17'b00010010101110001,
    17'b11101010010100100,
    17'b11110110101110001,
    17'b00001111010001111,
    17'b00001111000111101,
    17'b00000011100001010,
    17'b11111011100110011,
    17'b11110010000000000,
    17'b11110011010111000,
    17'b11111100101110001,
    17'b00100001110000101,
    17'b00110100000101001,
    17'b00100011110101110,
    17'b00011001000111101,
    17'b00001110000000000,
    17'b00100010111000011,
    17'b00100110010100100,
    17'b00101010011110110,
    17'b00101011100110011,
    17'b00101011111010111,
    17'b00110000000101001,
    17'b00101011100110011,
    17'b00101011110101110,
    17'b00101011011100001,
    17'b00101011000111101,
    17'b00101100000101001,
    17'b00101101011100001,
    17'b00101001110101110,
    17'b00100010111101100,
    17'b00011010011001101,
    17'b00010000010100100,
    17'b00001100101110001,
    17'b00001101100110011,
    17'b00010010001111011,
    17'b00011000111000011,
    17'b01001010101001000,
    17'b00110110010100100,
    17'b00110001110101110,
    17'b00110001101011100,
    17'b00101010101001000,
    17'b00101010101110001,
    17'b00101000101110001,
    17'b00101000001111011,
    17'b00101000011110110,
    17'b00101000011110110,
    17'b00101000011001101,
    17'b00101000101110001,
    17'b00101110001111011,
    17'b00110000011001101,
    17'b00101110100011111,
    17'b00101100011001101,
    17'b00100111001100110,
    17'b00100010111101100,
    17'b00011111111010111,
    17'b00011101100001010,
    17'b00011100011001101,
    17'b00011100110011010,
    17'b00011110000000000,
    17'b00011111100110011,
    17'b00110011101011100,
    17'b00101111100001010,
    17'b00101011010111000,
    17'b00101100001010010,
    17'b00101010011001101,
    17'b00101001100110011,
    17'b00101001001100110,
    17'b00101000101110001,
    17'b00101000001010010,
    17'b00101000000101001,
    17'b00101000000000000,
    17'b00100111110101110,
    17'b00101000110011010,
    17'b00101001011100001,
    17'b00101000011001101,
    17'b00101000000000000,
    17'b00100111010111000,
    17'b00100110000101001,
    17'b00100101010111000,
    17'b00100100011110110,
    17'b00100011010111000,
    17'b00100011000111101,
    17'b00100011100001010,
    17'b00101000111000011,
    17'b00101010101001000,
    17'b00101000011110110,
    17'b00101000110011010,
    17'b00100111010111000,
    17'b00100110101110001,
    17'b00100111100110011,
    17'b00100110011001101,
    17'b00100101000111101,
    17'b00100101110101110,
    17'b00100100111101100,
    17'b00100100010100100,
    17'b00101001110000101,
    17'b00101011000111101,
    17'b00101111010111000,
    17'b00101100011001101,
    17'b00111000110011010,
    17'b00011111100110011,
    17'b00101010011001101,
    17'b00100101110000101,
    17'b00011000010100100,
    17'b00001010001111011,
    17'b00001011001100110,
    17'b00111001010001111,
    17'b01001001111010111,
    17'b01011011100001010,
    17'b01001110101001000,
    17'b00110101000111101,
    17'b00101011111010111,
    17'b00110001001100110,
    17'b00111011001100110,
    17'b01000010001111011,
    17'b01000110000101001,
    17'b01001010101001000,
    17'b01001111000111101,
    17'b01001110000000000,
    17'b01000100110011010,
    17'b00110100111101100,
    17'b00100100000000000,
    17'b00011111000010100,
    17'b00011100111101100,
    17'b00011011100001010,
    17'b00011010101110001,
    17'b00011010101001000,
    17'b00011011011100001,
    17'b00011101100001010,
    17'b00100000110011010,
    17'b00100101011100001,
    17'b00101001010001111,
    17'b00101100101110001,
    17'b00110001110000101,
    17'b00110101101011100,
    17'b00111000100011111,
    17'b00111001000010100,
    17'b00111000011001101,
    17'b00110111100001010,
    17'b00110111010001111,
    17'b00110111110000101,
    17'b00111000010100100,
    17'b00110111110000101,
    17'b00110100000101001,
    17'b00101110101001000,
    17'b00101101100001010,
    17'b00110000111000011,
    17'b00110001011100001,
    17'b00110001110101110,
    17'b00110001110000101,
    17'b00110010011001101,
    17'b00110101000111101,
    17'b00110111110000101,
    17'b00111010110011010,
    17'b00111111010111000,
    17'b01000011000111101,
    17'b01000110011110110,
    17'b01000111110000101,
    17'b01000101110101110,
    17'b01000000111000011,
    17'b00111100111101100,
    17'b00111001111010111,
    17'b00111001110101110,
    17'b00111000111000011,
    17'b00111000001010010,
    17'b00110110110011010,
    17'b00110010100011111,
    17'b00101110001111011,
    17'b00101011100001010,
    17'b00101001100001010,
    17'b00100101010111000,
    17'b00001010100011111,
    17'b00000101110000101,
    17'b00001100001111011,
    17'b00100000011001101,
    17'b00101100011001101,
    17'b00110110111101100,
    17'b00111000011001101,
    17'b00110110011110110,
    17'b00111111010001111,
    17'b01001111011100001,
    17'b01010111011100001,
    17'b01010101010001111,
    17'b01011100001010010,
    17'b01010001011100001,
    17'b01000100001111011,
    17'b01000010001111011,
    17'b00100101101011100,
    17'b00110011000111101,
    17'b00111001011100001,
    17'b00110100101001000,
    17'b00101101011100001,
    17'b00100110000101001,
    17'b00011110101001000,
    17'b00010101100001010,
    17'b00001011010111000,
    17'b00000110001010010,
    17'b00000010111101100,
    17'b00000110101110001,
    17'b00001100001010010,
    17'b00000010110011010,
    17'b11110110010100100,
    17'b11101100011001101,
    17'b11100000001010010,
    17'b11010000110011010,
    17'b10111111000111101,
    17'b10110011100001010,
    17'b10110010001010010,
    17'b10110001100110011,
    17'b11100010110011010,
    17'b01110101010111000,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b00101101100110011,
    17'b11011101110101110,
    17'b11010101011100001,
    17'b11101010011001101,
    17'b00001010101110001,
    17'b00101101101011100,
    17'b01001010101001000,
    17'b01001011010111000,
    17'b01000100001010010,
    17'b00110111010001111,
    17'b00011101011100001,
    17'b00000111110000101,
    17'b11110101010001111,
    17'b11101000110011010,
    17'b11100001101011100,
    17'b11011100101110001,
    17'b11011111110101110,
    17'b11101000111000011,
    17'b11110110110011010,
    17'b00001000011110110,
    17'b00010001111010111,
    17'b00010101111010111,
    17'b00011001000111101,
    17'b00011010000101001,
    17'b00010001000010100,
    17'b00001010000000000,
    17'b00000100111101100,
    17'b00000000100011111,
    17'b11110111000010100,
    17'b11101100011110110,
    17'b11100000101110001,
    17'b11011000000101001,
    17'b11010100011110110,
    17'b11010110101110001,
    17'b11011000111101100,
    17'b11011010100011111,
    17'b11011011000111101,
    17'b11011001110000101,
    17'b11011000111000011,
    17'b11011000000101001,
    17'b11010110011001101,
    17'b11010100011001101,
    17'b11010100001111011,
    17'b11010101000010100,
    17'b11010111100001010,
    17'b11011001100110011,
    17'b11011010001111011,
    17'b11011000111101100,
    17'b11011000101110001,
    17'b11011010001010010,
    17'b11011100011001101,
    17'b11011101000111101,
    17'b11011110100011111,
    17'b11011101001100110,
    17'b11011011001100110,
    17'b11011000111000011,
    17'b11010101000111101,
    17'b11010001100001010,
    17'b11001010100011111,
    17'b11000100011110110,
    17'b10111100001111011,
    17'b10110100000101001,
    17'b10101101111010111,
    17'b10101110001010010,
    17'b10110010110011010,
    17'b10111010001111011,
    17'b11000001100110011,
    17'b11001000001111011,
    17'b11001001100001010,
    17'b11000111011100001,
    17'b11000010101110001,
    17'b10111010010100100,
    17'b10110100100011111,
    17'b10110000101110001,
    17'b10101110100011111,
    17'b10101110000000000,
    17'b10101111010111000,
    17'b10110010000101001,
    17'b10110110001111011,
    17'b10111011010001111,
    17'b11000010101001000,
    17'b11001000001111011,
    17'b11001110111000011,
    17'b11010100101110001,
    17'b11011001100001010,
    17'b11011101011100001,
    17'b11100000111101100,
    17'b11100110011110110,
    17'b11101010100011111,
    17'b11101111010001111,
    17'b11110011101011100,
    17'b11111101001100110,
    17'b00000010011001101,
    17'b00000011000010100,
    17'b00000001000111101,
    17'b11111000101001000,
    17'b11100011010001111,
    17'b10101111011100001,
    17'b10111000001111011,
    17'b11000110001111011,
    17'b11001100101110001,
    17'b11010010000101001,
    17'b11010010001010010,
    17'b11010100000101001,
    17'b11011011010111000,
    17'b11110111001100110,
    17'b11110111101011100,
    17'b11101100000000000,
    17'b11100101000111101,
    17'b11100001010111000,
    17'b11100000001111011,
    17'b11100000110011010,
    17'b11100001001100110,
    17'b11100010001010010,
    17'b11100011000010100,
    17'b11100011000010100,
    17'b11100011100001010,
    17'b11100100000000000,
    17'b11100110011110110,
    17'b11101001001100110,
    17'b11101010111101100,
    17'b11101101000111101,
    17'b11110100010100100,
    17'b11110111100110011,
    17'b11111010000000000,
    17'b11111101000111101,
    17'b11111111001100110,
    17'b11111110001010010,
    17'b11111110011001101,
    17'b00000001110101110,
    17'b00000011100001010,
    17'b00000101101011100,
    17'b00000101001100110,
    17'b00001000111101100,
    17'b00001000101001000,
    17'b00001011000111101,
    17'b00001100101110001,
    17'b00001110011001101,
    17'b00010000100011111,
    17'b00010010111000011,
    17'b00010011000010100,
    17'b00010100100011111,
    17'b00010100011001101,
    17'b00010101010111000,
    17'b00010100011001101,
    17'b00010010001010010,
    17'b00001111010111000,
    17'b00010101010111000,
    17'b00010110011001101,
    17'b00011010111101100,
    17'b00011110010100100,
    17'b00100010000101001,
    17'b00100100010100100,
    17'b00011101110101110,
    17'b00010101111010111,
    17'b00010001111010111,
    17'b00001110001010010,
    17'b00001011010111000,
    17'b00001010101001000,
    17'b00001101001100110,
    17'b00010010100011111,
    17'b00011010000000000,
    17'b00011110010100100,
    17'b00100000101001000,
    17'b00100010000101001,
    17'b00100010110011010,
    17'b00100010101110001,
    17'b00100011010001111,
    17'b00100011011100001,
    17'b00100100010100100,
    17'b00100110011110110,
    17'b00101000000101001,
    17'b00101010111000011,
    17'b00101100111101100,
    17'b00101101010001111,
    17'b00101100010100100,
    17'b00101010001111011,
    17'b00101001011100001,
    17'b00101011000010100,
    17'b00100010111000011,
    17'b00101010001010010,
    17'b00101110101110001,
    17'b00101011011100001,
    17'b00101011000111101,
    17'b00101011110101110,
    17'b00100111011100001,
    17'b00101001010001111,
    17'b00100110011001101,
    17'b00100011101011100,
    17'b00100010011001101,
    17'b00100000010100100,
    17'b00011110000101001,
    17'b00011010011001101,
    17'b00010111010111000,
    17'b00010100111101100,
    17'b00010010001111011,
    17'b00010000000101001,
    17'b00001110001010010,
    17'b00001101010001111,
    17'b00001011010111000,
    17'b00001011001100110,
    17'b00001010011001101,
    17'b00001001111010111,
    17'b00001011000010100,
    17'b00001010100011111,
    17'b00001000101001000,
    17'b00000110100011111,
    17'b00000011100001010,
    17'b00000001110101110,
    17'b00000000001010010,
    17'b11111110101001000,
    17'b11111110111101100,
    17'b11111110101001000,
    17'b11111110001010010,
    17'b11111110101001000,
    17'b11111111010001111,
    17'b00000000000101001,
    17'b00000001001100110,
    17'b00000001100001010,
    17'b00000001110101110,
    17'b00000001100110011,
    17'b00000001101011100,
    17'b00000010110011010,
    17'b00000011000010100,
    17'b00000011001100110,
    17'b00000011010001111,
    17'b00000010000000000,
    17'b00000010001111011,
    17'b00000010000000000,
    17'b00000000111101100,
    17'b00000000000000000,
    17'b11111111100001010,
    17'b11111111010001111,
    17'b11111110011001101,
    17'b11111110111000011,
    17'b11111111011100001,
    17'b00000000000000000,
    17'b00000001000010100,
    17'b00000010100011111,
    17'b00000100101001000,
    17'b00000101100110011,
    17'b00000101000111101,
    17'b00000111011100001,
    17'b00001011001100110,
    17'b00000100111000011,
    17'b00000101000010100,
    17'b00010010000000000,
    17'b00010101110101110,
    17'b00010001100110011,
    17'b00010000000000000,
    17'b00011001111010111,
    17'b00011010101001000,
    17'b00011000101001000,
    17'b00011110101001000,
    17'b00010101010001111,
    17'b00100000001010010,
    17'b00101000101001000,
    17'b00100110101110001,
    17'b00100011110000101,
    17'b00100000001111011,
    17'b00001111000111101,
    17'b00100000100011111,
    17'b00011101010001111,
    17'b00001101111010111,
    17'b00010111000010100,
    17'b00010111000010100,
    17'b00011101110000101,
    17'b00011100001010010,
    17'b00100010000101001,
    17'b00101010101110001,
    17'b00101110100011111,
    17'b00111001100110011,
    17'b01000110010100100,
    17'b01000001101011100,
    17'b00110010110011010,
    17'b00101010001111011,
    17'b00101001111010111,
    17'b00001011010001111,
    17'b11101001110101110,
    17'b11101100000000000,
    17'b00001000110011010,
    17'b01000000101001000,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111111111010111,
    17'b00111011110101110,
    17'b00110000111101100,
    17'b00100011110101110,
    17'b00000000010100100,
    17'b11101011100110011,
    17'b11100100110011010,
    17'b11111110000101001,
    17'b00011111001100110,
    17'b00111100110011010,
    17'b01001001101011100,
    17'b00111010001010010,
    17'b00110011110101110,
    17'b00110100000101001,
    17'b00111100100011111,
    17'b01011101111010111,
    17'b01001111010001111,
    17'b00111111010111000,
    17'b00111001001100110,
    17'b01001100100011111,
    17'b01101000000000000,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111110010100100,
    17'b01110100001010010,
    17'b01101110101110001,
    17'b01100001111010111,
    17'b00111010100011111,
    17'b00101011010111000,
    17'b00111100011001101,
    17'b01010011100110011,
    17'b01100101010001111,
    17'b01101110000000000,
    17'b01111000101001000,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01100011110101110,
    17'b01001001010111000,
    17'b00010001001100110,
    17'b11110100111101100,
    17'b11101000100011111,
    17'b11101010000101001,
    17'b11111001011100001,
    17'b00001101010111000,
    17'b00011100010100100,
    17'b00100101100110011,
    17'b00101111111010111,
    17'b00110110101001000,
    17'b00111000010100100,
    17'b01000000011110110,
    17'b01001001100110011,
    17'b01000010001111011,
    17'b00111000101110001,
    17'b00100101010111000,
    17'b00011111011100001,
    17'b00001110011001101,
    17'b00001101100001010,
    17'b00000101110101110,
    17'b00000100111000011,
    17'b00000001101011100,
    17'b11111101000111101,
    17'b00001000000000000,
    17'b00010100110011010,
    17'b00011000111000011,
    17'b00010111100110011,
    17'b00010011100110011,
    17'b00010001000010100,
    17'b00010000111101100,
    17'b00001011000010100,
    17'b00000001000010100,
    17'b11110111100110011,
    17'b11111010011001101,
    17'b11111000111101100,
    17'b11110100111101100,
    17'b11111100010100100,
    17'b00000010101110001,
    17'b00000101000010100,
    17'b00000110100011111,
    17'b00001000001111011,
    17'b00001000110011010,
    17'b00001000100011111,
    17'b00001001000111101,
    17'b00001011001100110,
    17'b00001110001010010,
    17'b00010001011100001,
    17'b00010001110000101,
    17'b00010000001010010,
    17'b00001101011100001,
    17'b00001010000000000,
    17'b00000111100110011,
    17'b00000101010001111,
    17'b00000011001100110,
    17'b00000000000000000,
    17'b11111100101110001,
    17'b11111000010100100,
    17'b11110110011110110,
    17'b11101101011100001,
    17'b11100011111010111,
    17'b11100100111000011,
    17'b11100001001100110,
    17'b11011101010111000,
    17'b11011001110101110,
    17'b11010101111010111,
    17'b11001110001111011,
    17'b11001011010111000,
    17'b11001111010001111,
    17'b11001010101110001,
    17'b11001000001010010,
    17'b11000111110101110,
    17'b11001001101011100,
    17'b11001100111000011,
    17'b11010001111010111,
    17'b11010011011100001,
    17'b11010101110101110,
    17'b11010111111010111,
    17'b11001101011100001,
    17'b11010011100110011,
    17'b11010101001100110,
    17'b11010011000010100,
    17'b11011010101001000,
    17'b11010111100001010,
    17'b11001111100110011,
    17'b11001000101110001,
    17'b11010100101001000,
    17'b11001011110000101,
    17'b11010000001111011,
    17'b11001110101001000,
    17'b11010100110011010,
    17'b11000111010001111,
    17'b11011100000000000,
    17'b11011000101001000,
    17'b11011001110000101,
    17'b11011111101011100,
    17'b11100100010100100,
    17'b11101001000010100,
    17'b11101111100110011,
    17'b11110011101011100,
    17'b11110011110000101,
    17'b11110010001111011,
    17'b11101111100110011,
    17'b11101111011100001,
    17'b11101101100001010,
    17'b11101110000000000,
    17'b11101101100110011,
    17'b11101011110101110,
    17'b11101110110011010,
    17'b11101111110000101,
    17'b11101100000000000,
    17'b11101010101110001,
    17'b11101101110101110,
    17'b11110110101001000,
    17'b11111110101001000,
    17'b00000110001010010,
    17'b00001101000111101,
    17'b00010001000111101,
    17'b00010001001100110,
    17'b00010010000101001,
    17'b00010010000101001,
    17'b00010010001010010,
    17'b00010010011001101,
    17'b00010100011110110,
    17'b00010110111000011,
    17'b00011001001100110,
    17'b00011010001111011,
    17'b00011001000010100,
    17'b00011000011110110,
    17'b00010110101110001,
    17'b00010100100011111,
    17'b00010001111010111,
    17'b00001110101001000,
    17'b00010000001111011,
    17'b00010001100110011,
    17'b11110111110101110,
    17'b11101100001010010,
    17'b00001111100001010,
    17'b00100001000010100,
    17'b00100010001010010,
    17'b00100110001010010,
    17'b00110101010001111,
    17'b00111010110011010,
    17'b00111010011001101,
    17'b00111000100011111,
    17'b00110111010111000,
    17'b00111000000101001,
    17'b00111000000000000,
    17'b00110100100011111,
    17'b00101110000101001,
    17'b00111010000000000,
    17'b01000010100011111,
    17'b01001000111000011,
    17'b01011001001100110,
    17'b01011101010001111,
    17'b01010100111101100,
    17'b01010101010001111,
    17'b01011110000101001,
    17'b01100111110101110,
    17'b01101001101011100,
    17'b01100100001111011,
    17'b01011001000111101,
    17'b01010010001111011,
    17'b01000110001010010,
    17'b01000001010001111,
    17'b01010011010111000,
    17'b01011001110000101,
    17'b01100000011110110,
    17'b01100001100001010,
    17'b01011100010100100,
    17'b01010001010001111,
    17'b01001100011110110,
    17'b01001010101001000,
    17'b01001001110000101,
    17'b01001001101011100,
    17'b01001001100001010,
    17'b01000111111010111,
    17'b01000100111101100,
    17'b01000011000111101,
    17'b01000011000010100,
    17'b01000001100001010,
    17'b00111111010111000,
    17'b00111110000000000,
    17'b00111110011110110,
    17'b00111101111010111,
    17'b00111110110011010,
    17'b00111100000101001,
    17'b00110001100110011,
    17'b00101001110101110,
    17'b00100111001100110,
    17'b00101010001111011,
    17'b00110110000000000,
    17'b00111011100001010,
    17'b00111010100011111,
    17'b00110100110011010,
    17'b00101010001010010,
    17'b00100110000101001,
    17'b00101001000111101,
    17'b00101000110011010,
    17'b00100111010111000,
    17'b00100111110101110,
    17'b00101001001100110,
    17'b00101010101110001,
    17'b00101010011110110,
    17'b00101100011001101,
    17'b00110010111000011,
    17'b00111100111000011,
    17'b01001001111010111,
    17'b01001111111010111,
    17'b01001111110101110,
    17'b01001001001100110,
    17'b00100011010111000,
    17'b00100100100011111,
    17'b00101000010100100,
    17'b00110100111101100,
    17'b01000101110000101,
    17'b01010111001100110,
    17'b01100101101011100,
    17'b01101010101110001,
    17'b01100110110011010,
    17'b01010101111010111,
    17'b01000100110011010,
    17'b00110100011001101,
    17'b00100111000111101,
    17'b00100010011110110,
    17'b00100100111000011,
    17'b00101001100110011,
    17'b00101001110101110,
    17'b00100001100110011,
    17'b00001110001111011,
    17'b00000001100110011,
    17'b11111000100011111,
    17'b11110101110101110,
    17'b11111101110000101,
    17'b00001101010001111,
    17'b00011111000010100,
    17'b00110001000010100,
    17'b00111000001010010,
    17'b00111011010001111,
    17'b00111010011110110,
    17'b00111001011100001,
    17'b01001111110000101,
    17'b01101101010001111,
    17'b01111000110011010,
    17'b01101000010100100,
    17'b01010110000000000,
    17'b01000011110101110,
    17'b00110001111010111,
    17'b01010111011100001,
    17'b01110010110011010,
    17'b01010111101011100,
    17'b00110111000010100,
    17'b00100001000010100,
    17'b00010111100001010,
    17'b00010000111000011,
    17'b00010100110011010,
    17'b00100110110011010,
    17'b00110010010100100,
    17'b00110111000010100,
    17'b00110111010001111,
    17'b00110101000111101,
    17'b00110100001010010,
    17'b00110011100001010,
    17'b00110010001010010,
    17'b00110011110101110,
    17'b00111000011001101,
    17'b00110111001100110,
    17'b00101110101001000,
    17'b00100010100011111,
    17'b00100000000101001,
    17'b00100010011001101,
    17'b00100101010001111,
    17'b00100111100001010,
    17'b00100111001100110,
    17'b00100100011001101,
    17'b00011111110000101,
    17'b00011010001010010,
    17'b00010011010111000,
    17'b00001111110000101,
    17'b00001101100110011,
    17'b00001100011001101,
    17'b00001100001111011,
    17'b00001100100011111,
    17'b00001100101110001,
    17'b00001100101001000,
    17'b00001100001010010,
    17'b00001011111010111,
    17'b00001101000010100,
    17'b00001110110011010,
    17'b00010000011001101,
    17'b00010001111010111,
    17'b00010010000000000,
    17'b00010000101110001,
    17'b00001110111101100,
    17'b00001101000111101,
    17'b00001101000010100,
    17'b00001110111101100,
    17'b00010001000010100,
    17'b00010010001111011,
    17'b00010001000010100,
    17'b00001101100001010,
    17'b00001000000000000,
    17'b00000010000000000,
    17'b11111010111101100,
    17'b11110111010111000,
    17'b11110100101110001,
    17'b11110010110011010,
    17'b11110001000111101,
    17'b11110010001010010,
    17'b11110000011110110,
    17'b11100111100001010,
    17'b11100110010100100,
    17'b11101001000010100,
    17'b11101011011100001,
    17'b11101110000101001,
    17'b11101110111101100,
    17'b11110000111101100,
    17'b11110100001111011,
    17'b11111000101001000,
    17'b11111010101110001,
    17'b11111011000010100,
    17'b11111001010111000,
    17'b11110101010001111,
    17'b11110001001100110,
    17'b11101100011110110,
    17'b11100111000111101,
    17'b11100000011110110,
    17'b11011100100011111,
    17'b11011011000010100,
    17'b11011011110101110,
    17'b11011011100110011,
    17'b11011001011100001,
    17'b11010110110011010,
    17'b11010011110000101,
    17'b11010000001111011,
    17'b11001101110000101,
    17'b11000111001100110,
    17'b10111011011100001,
    17'b10101110111101100,
    17'b10110000101001000,
    17'b10111010001111011,
    17'b11000011101011100,
    17'b11001000011001101,
    17'b11001000011110110,
    17'b11000101110000101,
    17'b11000001100110011,
    17'b10111100001111011,
    17'b10110101110000101,
    17'b10110010101110001,
    17'b10110001000111101,
    17'b10101111110101110,
    17'b10101110011001101,
    17'b10101101010111000,
    17'b10101101111010111,
    17'b10110001000010100,
    17'b10110100010100100,
    17'b10110111000111101,
    17'b10110111111010111,
    17'b10110110000101001,
    17'b10110010101001000,
    17'b10110001001100110,
    17'b10110001010111000,
    17'b10110010101001000,
    17'b10110100110011010,
    17'b10110111000111101,
    17'b10111010011001101,
    17'b10111100011110110,
    17'b10111101100001010,
    17'b10111110000101001,
    17'b10111110000101001,
    17'b10111101101011100,
    17'b10111101101011100,
    17'b10111101110000101,
    17'b10111101110000101,
    17'b10111110001010010,
    17'b10111111010111000,
    17'b11000011010111000,
    17'b11000110101001000,
    17'b11001011000010100,
    17'b11010000111000011,
    17'b11010101100110011,
    17'b11011010011001101,
    17'b11011101010001111,
    17'b11011110000101001,
    17'b11011101110101110,
    17'b11011011110000101,
    17'b11011011000010100,
    17'b11011010101110001,
    17'b11011011000010100,
    17'b11011010000000000,
    17'b11011011010001111,
    17'b11011101111010111,
    17'b11011110010100100,
    17'b11011011001100110,
    17'b11011100010100100,
    17'b11100100001010010,
    17'b11101111100110011,
    17'b11111010111101100,
    17'b00000010101001000,
    17'b00000101110000101,
    17'b00001000000000000,
    17'b00001001010111000,
    17'b00001011000111101,
    17'b00001100011110110,
    17'b00000100111000011,
    17'b00000000000101001,
    17'b11111100111101100,
    17'b11111010001010010,
    17'b11111001010001111,
    17'b11111010011001101,
    17'b11111100001111011,
    17'b11111110101110001,
    17'b00000001111010111,
    17'b00000011010111000,
    17'b00000011110000101,
    17'b00000010111101100,
    17'b00000000101001000,
    17'b11100110000000000,
    17'b11001111000111101,
    17'b11100001111010111,
    17'b11111010111101100,
    17'b00010000111000011,
    17'b00100101000111101,
    17'b00010100001111011,
    17'b00010010001111011,
    17'b00011001000111101,
    17'b00100010110011010,
    17'b00101110110011010,
    17'b00110000010100100,
    17'b00101111001100110,
    17'b00101011110000101,
    17'b00101011010111000,
    17'b00101100011110110,
    17'b00101111110101110,
    17'b00110100001111011,
    17'b00110011000111101,
    17'b00110010011110110,
    17'b00110011010001111,
    17'b00110010101110001,
    17'b00110010110011010,
    17'b00110011110101110,
    17'b00110011100001010,
    17'b00110010011110110,
    17'b00110000111000011,
    17'b00101110111101100,
    17'b00101100001010010,
    17'b00101010001010010,
    17'b00100111000010100,
    17'b00100100011001101,
    17'b00100011100110011,
    17'b00100001110101110,
    17'b00010011101011100,
    17'b00010001111010111,
    17'b00010011110101110,
    17'b00100100101110001,
    17'b00110111110101110,
    17'b01001100011001101,
    17'b01010101011100001,
    17'b01010011111010111,
    17'b01000110100011111,
    17'b00110101011100001,
    17'b00100111100001010,
    17'b00011001100110011,
    17'b00010011010001111,
    17'b00011110101001000,
    17'b00101101101011100,
    17'b01000010010100100,
    17'b01010111100001010,
    17'b01100111100001010,
    17'b01101110000000000,
    17'b01100110001010010,
    17'b01011000000000000,
    17'b01001000000101001,
    17'b00111001010111000,
    17'b00101010111000011,
    17'b00100100011001101,
    17'b00100000111000011,
    17'b00011111010001111,
    17'b00011111010111000,
    17'b00100000111101100,
    17'b00100010101001000,
    17'b00100011110101110,
    17'b00100100101110001,
    17'b00100100111101100,
    17'b00100101100110011,
    17'b00100110100011111,
    17'b00100111111010111,
    17'b00101001001100110,
    17'b00101010101001000,
    17'b00101100101001000,
    17'b00101110000101001,
    17'b00101111011100001,
    17'b00110000110011010,
    17'b00110010101001000,
    17'b00110101110000101,
    17'b00111000011001101,
    17'b00111010001010010,
    17'b00111010111101100,
    17'b00111010001111011,
    17'b00111000111101100,
    17'b00110111111010111,
    17'b00110111110000101,
    17'b00110111110000101,
    17'b00110111000111101,
    17'b00110101100110011,
    17'b00110011100110011,
    17'b00110001010001111,
    17'b00101110101001000,
    17'b00101101100001010,
    17'b00101110000101001,
    17'b00101111101011100,
    17'b00110010001111011,
    17'b00110110011110110,
    17'b00111000011110110,
    17'b00111010001111011,
    17'b00111001011100001,
    17'b00111000111101100,
    17'b00111001100001010,
    17'b00111100100011111,
    17'b01000000111101100,
    17'b01000011001100110,
    17'b01000101001100110,
    17'b01000110000101001,
    17'b01000100100011111,
    17'b01000010010100100,
    17'b01000010111000011,
    17'b01000010010100100,
    17'b01000001111010111,
    17'b01000011100001010,
    17'b01000100111101100,
    17'b01000110000101001,
    17'b01000110001111011,
    17'b01000101101011100,
    17'b01000011101011100,
    17'b01000010111101100,
    17'b01000000101001000,
    17'b00111110011001101,
    17'b00111011011100001,
    17'b00111011010001111,
    17'b00111011000111101,
    17'b00111011010001111,
    17'b00111101110000101,
    17'b01000000000000000,
    17'b01000010100011111,
    17'b01000101000111101,
    17'b01000110001111011,
    17'b01000101111010111,
    17'b01000110100011111,
    17'b01000101100110011,
    17'b01000100110011010,
    17'b01000100101110001,
    17'b01000100001111011,
    17'b01000011000111101,
    17'b01000001100110011,
    17'b01000000001111011,
    17'b00111111000010100,
    17'b00111101001100110,
    17'b00111011010001111,
    17'b00111000100011111,
    17'b00110100110011010,
    17'b00110000011110110,
    17'b00101010101110001,
    17'b00100110110011010,
    17'b00100011101011100,
    17'b00100001111010111,
    17'b00100001101011100,
    17'b00100011010111000,
    17'b00100110001010010,
    17'b00101010001111011,
    17'b00101111000010100,
    17'b00110100101110001,
    17'b00111001011100001,
    17'b00111100000000000,
    17'b00111100101110001,
    17'b00111110111000011,
    17'b00111110111101100,
    17'b00111110011001101,
    17'b00111110010100100,
    17'b00111100110011010,
    17'b00111010111101100,
    17'b00110111111010111,
    17'b00110101010001111,
    17'b00110010111000011,
    17'b00101111110101110,
    17'b00101100001111011,
    17'b00101000000000000,
    17'b00101011110000101,
    17'b00110111110000101,
    17'b00111111101011100,
    17'b01000010001010010,
    17'b01000001000111101,
    17'b00111111101011100,
    17'b00111101001100110,
    17'b00110111001100110,
    17'b00110001111010111,
    17'b00101110001010010,
    17'b00101101000111101,
    17'b00101110011110110,
    17'b00110001111010111,
    17'b00110101100001010,
    17'b00111001110101110,
    17'b00111101101011100,
    17'b01000001000111101,
    17'b01000010011001101,
    17'b01000010100011111,
    17'b01000000111000011,
    17'b01000011111010111,
    17'b01000100110011010,
    17'b01000010001010010,
    17'b00111110100011111,
    17'b00111110101001000,
    17'b01000101010001111,
    17'b01001100011110110,
    17'b01010011110000101,
    17'b01011001001100110,
    17'b01011011110101110,
    17'b01011010011110110,
    17'b01010110011110110,
    17'b01001111011100001,
    17'b01001000101110001,
    17'b01000010011110110,
    17'b00111110001111011,
    17'b00111100000101001,
    17'b00111000111101100,
    17'b00110011100110011,
    17'b00110001011100001,
    17'b00110001110101110,
    17'b00110011000111101,
    17'b00110100111101100,
    17'b00110101000010100,
    17'b00110101000010100,
    17'b00110101001100110,
    17'b00110100000000000,
    17'b00101111100001010,
    17'b00101011101011100,
    17'b00101000001010010,
    17'b00100101000111101,
    17'b00100001010111000,
    17'b00011111001100110,
    17'b00011101100001010,
    17'b00011100011001101,
    17'b00011010001111011,
    17'b00011010010100100,
    17'b00011100101110001,
    17'b00100001010001111,
    17'b00100111111010111,
    17'b00110001000111101,
    17'b00110111011100001,
    17'b00111011101011100,
    17'b00111101101011100,
    17'b00111101000010100,
    17'b00111010110011010,
    17'b00110111001100110,
    17'b00110001110000101,
    17'b00101011001100110,
    17'b00100010000101001,
    17'b00011011110000101,
    17'b00010110011110110,
    17'b00010010111101100,
    17'b00010000011110110,
    17'b00001111110101110,
    17'b00001111010111000,
    17'b00001111010111000,
    17'b00001111110000101,
    17'b00010001110000101,
    17'b00010100000000000,
    17'b00010110111000011,
    17'b00011010001010010,
    17'b00011100110011010,
    17'b00011111110000101,
    17'b00100001100001010,
    17'b00100110011001101,
    17'b00110100001111011,
    17'b01001011010001111,
    17'b01101001101011100,
    17'b01110101101011100,
    17'b01110111100001010,
    17'b01110001000111101,
    17'b01100100011110110,
    17'b01001010101001000,
    17'b00110010110011010,
    17'b00011010111000011,
    17'b00000110111000011,
    17'b11110111011100001,
    17'b11110100100011111,
    17'b11110111000111101,
    17'b11111100111000011,
    17'b00000011110101110,
    17'b00001100100011111,
    17'b00010010110011010,
    17'b00011001001100110,
    17'b00011111110101110,
    17'b00100011010111000,
    17'b00100100000101001,
    17'b00011011000111101,
    17'b00000111110101110,
    17'b11110011000010100,
    17'b11101111101011100,
    17'b00000100000101001,
    17'b00011000101110001,
    17'b00101001010111000,
    17'b00110100010100100,
    17'b00110110101110001,
    17'b00101111000111101,
    17'b00100100101110001,
    17'b00011010010100100,
    17'b00010010101001000,
    17'b00010000000000000,
    17'b00010111000111101,
    17'b00011111101011100,
    17'b00101000000101001,
    17'b00101110001111011,
    17'b00110000111000011,
    17'b00101111010001111,
    17'b00101000000000000,
    17'b00100011110000101,
    17'b00100011101011100,
    17'b00100110010100100,
    17'b00100110101001000,
    17'b00100011100001010,
    17'b00011110110011010,
    17'b00011010000000000,
    17'b00011000101001000,
    17'b00011000010100100,
    17'b00010111101011100,
    17'b00010110011001101,
    17'b00010100001010010,
    17'b00001111010111000,
    17'b00001010011001101,
    17'b00000110111101100,
    17'b00000100011001101,
    17'b00000010101110001,
    17'b00000000111101100,
    17'b11111111000111101,
    17'b11111111010001111,
    17'b00000001001100110,
    17'b00000100001111011,
    17'b00000010100011111,
    17'b11111111001100110,
    17'b11111100010100100,
    17'b00000001100001010,
    17'b00000000011110110,
    17'b11111001010001111,
    17'b11101111001100110,
    17'b11101011110000101,
    17'b11101100111000011,
    17'b11110001000111101,
    17'b11110111000010100,
    17'b11111011010111000,
    17'b00000001001100110,
    17'b00001000111000011,
    17'b00010011000111101,
    17'b00011001001100110,
    17'b00011110000000000,
    17'b00100001010111000,
    17'b00100010011001101,
    17'b00011111110000101,
    17'b00011011100001010,
    17'b00011000000000000,
    17'b00010011000111101,
    17'b00001100001111011,
    17'b00001011000111101,
    17'b00001000011001101,
    17'b00000010100011111,
    17'b11111111100001010,
    17'b11111001100001010,
    17'b11111100001010010,
    17'b00000011110101110,
    17'b00001110000000000,
    17'b00011000011110110,
    17'b00011111000111101,
    17'b00101011001100110,
    17'b00110011101011100,
    17'b00111100101110001,
    17'b01000000101001000,
    17'b01000011010001111,
    17'b01000100111101100,
    17'b01000100100011111,
    17'b01000010010100100,
    17'b00111101101011100,
    17'b00111010111101100,
    17'b00111111110000101,
    17'b01001001000010100,
    17'b01010001100110011,
    17'b01010100001111011,
    17'b01010010110011010,
    17'b01001111100110011,
    17'b01001010101110001,
    17'b01001000011001101,
    17'b01000011100001010,
    17'b01000001000111101,
    17'b00110101110101110,
    17'b00101011100001010,
    17'b00100011110101110,
    17'b00011100010100100,
    17'b00010110001111011,
    17'b00011000100011111,
    17'b00011111011100001,
    17'b00100101010111000,
    17'b00101000001010010,
    17'b00100110111101100,
    17'b00100110000000000,
    17'b00101000011001101,
    17'b00101101011100001,
    17'b00101111011100001,
    17'b00101110111101100,
    17'b00101101110101110,
    17'b00101101011100001,
    17'b00101110100011111,
    17'b00110000110011010,
    17'b00110111111010111,
    17'b00111000100011111,
    17'b00110111100001010,
    17'b00110101100110011,
    17'b00110011110000101,
    17'b00110011000111101,
    17'b00110010110011010,
    17'b00110010101001000,
    17'b00110011010111000,
    17'b00110100011001101,
    17'b00110101101011100,
    17'b00110111000111101,
    17'b00111001001100110,
    17'b00111010111000011,
    17'b00111011011100001,
    17'b00111001100001010,
    17'b00110101100001010,
    17'b00101110101001000,
    17'b00100100111000011,
    17'b00011011000111101,
    17'b00011000111000011,
    17'b00011001010111000,
    17'b00011010010100100,
    17'b00011001000111101,
    17'b00010111111010111,
    17'b00010110110011010,
    17'b00010111000010100,
    17'b00010111101011100,
    17'b00010101111010111,
    17'b00010011000111101,
    17'b00001110011001101,
    17'b00000110001111011,
    17'b11111011100110011,
    17'b11110011011100001,
    17'b11110000101001000,
    17'b11110011111010111,
    17'b11111100000101001,
    17'b00000111000010100,
    17'b00010010101001000,
    17'b00011000110011010,
    17'b00011110110011010,
    17'b00100100001111011,
    17'b00101000101110001,
    17'b00101000011110110,
    17'b00100100111101100,
    17'b00011111000010100,
    17'b00011000100011111,
    17'b00010110100011111,
    17'b00010110000000000,
    17'b00010100110011010,
    17'b00010000111000011,
    17'b00001100111000011,
    17'b00001000100011111,
    17'b00000011010001111,
    17'b11111011111010111,
    17'b11110111000010100,
    17'b11110010101110001,
    17'b11101101001100110,
    17'b11101010000000000,
    17'b11101000000101001,
    17'b11101000000101001,
    17'b11101000000000000,
    17'b11101000011110110,
    17'b11101000111000011,
    17'b11101000111000011,
    17'b11101010010100100,
    17'b11101101111010111,
    17'b11101100111101100,
    17'b11101100010100100,
    17'b11101101010111000,
    17'b11101111000010100,
    17'b11110000101001000,
    17'b11110010011001101,
    17'b11110010010100100,
    17'b11110001001100110,
    17'b11101111000010100,
    17'b11101001110101110,
    17'b11100101001100110,
    17'b11100000111000011,
    17'b11011100100011111,
    17'b11011011001100110,
    17'b11011100000000000,
    17'b11011110000000000,
    17'b11011111110000101,
    17'b11011111000010100,
    17'b11011101010001111,
    17'b11011010111101100,
    17'b11010111111010111,
    17'b11010100000000000,
    17'b11010001110101110,
    17'b11010000011110110,
    17'b11001111000010100,
    17'b11001100110011010,
    17'b11001010101110001,
    17'b11001001100001010,
    17'b11001001111010111,
    17'b11001101101011100,
    17'b11010001110000101,
    17'b11010100101110001,
    17'b11010101011100001,
    17'b11010100101001000,
    17'b11010101000111101,
    17'b11010110110011010,
    17'b11010111110101110,
    17'b11010111100001010,
    17'b11010110000101001,
    17'b11010011100001010,
    17'b11010000100011111,
    17'b11001110010100100,
    17'b11001101110000101,
    17'b11001101011100001,
    17'b11001100111101100,
    17'b11001100000000000,
    17'b11001010111101100,
    17'b11001001101011100,
    17'b11000111110101110,
    17'b11000110001010010,
    17'b11000100101001000,
    17'b11000011111010111,
    17'b11000101111010111,
    17'b11000110111000011,
    17'b11000111100001010,
    17'b11000111110101110,
    17'b11000111110101110,
    17'b11000111001100110,
    17'b11000110010100100,
    17'b11000101010001111,
    17'b11000100100011111,
    17'b11000100000101001,
    17'b11000011111010111,
    17'b11000011110000101,
    17'b11000100010100100,
    17'b11000100111000011,
    17'b11000101000010100,
    17'b11000100101110001,
    17'b11000100001111011,
    17'b11000100000000000,
    17'b11000011110101110,
    17'b11000011100110011,
    17'b11000101001100110,
    17'b11001011010111000,
    17'b11011010000000000,
    17'b11011100011001101,
    17'b11010101010001111,
    17'b11001111000111101,
    17'b11001100000101001,
    17'b11001110001010010,
    17'b11010001010001111,
    17'b11010011010111000,
    17'b11010101111010111,
    17'b11011010110011010,
    17'b11011110000000000,
    17'b11011111100001010,
    17'b11100000101110001,
    17'b11100001110000101,
    17'b11100010100011111,
    17'b11100011001100110,
    17'b11100001111010111,
    17'b11011110110011010,
    17'b11011100111000011,
    17'b11011111011100001,
    17'b11100000101001000,
    17'b11100001110101110,
    17'b11100100011110110,
    17'b11100101100110011,
    17'b11100100011001101,
    17'b11100100111000011,
    17'b11100011110101110,
    17'b11011011101011100,
    17'b11011000101110001,
    17'b11010101111010111,
    17'b11011011000111101,
    17'b11001100011110110,
    17'b11001001000010100,
    17'b11010000111101100,
    17'b11000011100110011,
    17'b10101100111101100,
    17'b10001101011100001,
    17'b10111100111000011,
    17'b11110000100011111,
    17'b00001000001010010,
    17'b00000111100001010,
    17'b00000010101110001,
    17'b00000011000010100,
    17'b00001010000000000,
    17'b00010010111101100,
    17'b00011010011001101,
    17'b00011111010111000,
    17'b00100010111101100,
    17'b00100100101110001,
    17'b00100011010111000,
    17'b00100000010100100,
    17'b00011110101110001,
    17'b00011100010100100,
    17'b00011001100001010,
    17'b00010110111101100,
    17'b00010100101001000,
    17'b00010010000101001,
    17'b00010000001010010,
    17'b00001110011001101,
    17'b00001100101001000,
    17'b00001011100001010,
    17'b00001011010001111,
    17'b11111001100001010,
    17'b11011000011110110,
    17'b11011000111101100,
    17'b11111111100110011,
    17'b00101001110000101,
    17'b00101100010100100,
    17'b00100011111010111,
    17'b00100000101110001,
    17'b00101000010100100,
    17'b00101101010001111,
    17'b00101011110101110,
    17'b00100111011100001,
    17'b00100101110101110,
    17'b00101001101011100,
    17'b00101101000111101,
    17'b00110011110000101,
    17'b00111110011110110,
    17'b00111111010001111,
    17'b00111011011100001,
    17'b00110100110011010,
    17'b00101000110011010,
    17'b00011111010111000,
    17'b00010110101110001,
    17'b00001010101110001,
    17'b00000110110011010,
    17'b11111110101110001,
    17'b11111011100001010,
    17'b00000000100011111,
    17'b00001001110101110,
    17'b00001000000101001,
    17'b00000001010001111,
    17'b11111101000010100,
    17'b11111100101110001,
    17'b11111011110000101,
    17'b11111110100011111,
    17'b00001010111101100,
    17'b00010010110011010,
    17'b00010100001111011,
    17'b00010000111101100,
    17'b00010110111000011,
    17'b00010111000111101,
    17'b00001011010111000,
    17'b11111111011100001,
    17'b11110010111000011,
    17'b11100011111010111,
    17'b11100010101001000,
    17'b11100110110011010,
    17'b11100101001100110,
    17'b11101010101110001,
    17'b11101000110011010,
    17'b11100111100001010,
    17'b11100101001100110,
    17'b11100010100011111,
    17'b11011111101011100,
    17'b11011100010100100,
    17'b11011001110101110,
    17'b11010111001100110,
    17'b11010100000101001,
    17'b11001110111101100,
    17'b11001010101110001,
    17'b11000110001010010,
    17'b11000010100011111,
    17'b10111110111101100,
    17'b10111100111000011,
    17'b10111011100001010,
    17'b10111010100011111,
    17'b10111010101110001,
    17'b10111011101011100,
    17'b10111100010100100,
    17'b10111100010100100,
    17'b10111100011001101,
    17'b10111100001111011,
    17'b10111100000101001,
    17'b10111011000111101,
    17'b10111010001111011,
    17'b10111010000101001,
    17'b10111001110101110,
    17'b10110111111010111,
    17'b10111000110011010,
    17'b10111010000101001,
    17'b10111001010111000,
    17'b10110110001010010,
    17'b10110110101001000,
    17'b10110110101001000,
    17'b10110110110011010,
    17'b10111000000101001,
    17'b10111000011001101,
    17'b10110111000111101,
    17'b10110111010111000,
    17'b10110111000010100,
    17'b10110110111000011,
    17'b10110110110011010,
    17'b10110100000101001,
    17'b10110010011001101,
    17'b10110010111101100,
    17'b10101110101110001,
    17'b10101010011001101,
    17'b10101101000111101,
    17'b10101110111101100,
    17'b10101101100110011,
    17'b10101100110011010,
    17'b10101111010001111,
    17'b10110010100011111,
    17'b10110100101110001,
    17'b10110111010111000,
    17'b10111000011001101,
    17'b10111001010001111,
    17'b10110110000000000,
    17'b10110100001111011,
    17'b10110101110101110,
    17'b10110101010001111,
    17'b10110100111000011,
    17'b10011110111000011,
    17'b10011000110011010,
    17'b10000000000000000,
    17'b10000000000000000,
    17'b10000000000000000,
    17'b10000111000111101,
    17'b10001011100001010,
    17'b10001101000111101,
    17'b10000100101110001,
    17'b10010111100001010,
    17'b10010111110000101,
    17'b10011110101110001,
    17'b10101011110101110,
    17'b10110011100001010,
    17'b10110001010001111,
    17'b10110101100001010,
    17'b10111101011100001,
    17'b11000100101110001,
    17'b11001001110000101,
    17'b11001000110011010,
    17'b11000111001100110,
    17'b11000110011110110,
    17'b11000111100001010,
    17'b11001010000000000,
    17'b11001011110101110,
    17'b11001100101110001,
    17'b11001101101011100,
    17'b11001111110101110,
    17'b11010010001010010,
    17'b11010001100110011,
    17'b11001101001100110,
    17'b11001110000000000,
    17'b11010001100001010,
    17'b11010010101110001,
    17'b11010010011001101,
    17'b11010100010100100,
    17'b11011100101001000,
    17'b11100000101110001,
    17'b11011110101110001,
    17'b11011011110101110,
    17'b11011000101001000,
    17'b11100000110011010,
    17'b11100001100001010,
    17'b11011101001100110,
    17'b11011101010001111,
    17'b11011001011100001,
    17'b11011100011001101,
    17'b11011101100001010,
    17'b11100000010100100,
    17'b11100010111000011,
    17'b11100000000101001,
    17'b11011100011110110,
    17'b11100001001100110,
    17'b11100011110000101,
    17'b11100100000000000,
    17'b11100110110011010,
    17'b11101100010100100,
    17'b11110001110101110,
    17'b11110100101110001,
    17'b11111000101110001,
    17'b11111110001111011,
    17'b00000101001100110,
    17'b00001110100011111,
    17'b00011000111101100,
    17'b00011100011110110,
    17'b00010011110000101,
    17'b00000111010001111,
    17'b11111111111010111,
    17'b11111111011100001,
    17'b00001001111010111,
    17'b00010100111000011,
    17'b00010011000010100,
    17'b00010001101011100,
    17'b00010010101110001,
    17'b00010101011100001,
    17'b00010110101110001,
    17'b00010111001100110,
    17'b00100101010111000,
    17'b01111111111111111,
    17'b01110000111000011,
    17'b01000101101011100,
    17'b00111000011110110,
    17'b00101110001111011,
    17'b00100110111000011,
    17'b00100001110101110,
    17'b00011110110011010,
    17'b00100101000111101,
    17'b00011111001100110,
    17'b00011011001100110,
    17'b00010110100011111,
    17'b00010111011100001,
    17'b00010101001100110,
    17'b00001000110011010,
    17'b00000001110101110,
    17'b00000101100110011,
    17'b00001100110011010,
    17'b00010000111000011,
    17'b00010100001010010,
    17'b00010110011110110,
    17'b00010111010111000,
    17'b00010110000000000,
    17'b00010110101110001,
    17'b00010110001010010,
    17'b00001111110101110,
    17'b00001001100110011,
    17'b00000100111101100,
    17'b00000010000101001,
    17'b00000001001100110,
    17'b00000001010001111,
    17'b00000010111101100,
    17'b00000101010001111,
    17'b00000111111010111,
    17'b00001010010100100,
    17'b00001010110011010,
    17'b00001010001111011,
    17'b00000110000101001,
    17'b00000110110011010,
    17'b00000111100110011,
    17'b00001010010100100,
    17'b00010000101001000,
    17'b00010110000101001,
    17'b00010111101011100,
    17'b00011010111101100,
    17'b00011011110000101,
    17'b00011001000010100,
    17'b00010100100011111,
    17'b00010000011110110,
    17'b00010000011001101,
    17'b00010001000010100,
    17'b00010001110000101,
    17'b00010001111010111,
    17'b00010000100011111,
    17'b00001110010100100,
    17'b00001100111101100,
    17'b00001011010001111,
    17'b00001100001010010,
    17'b00010001000010100,
    17'b00011001001100110,
    17'b00011101001100110,
    17'b00011111111010111,
    17'b00100001000010100,
    17'b00100001000111101,
    17'b00100000011001101,
    17'b00011111110000101,
    17'b00011101111010111,
    17'b00011011010001111,
    17'b00011000000000000,
    17'b00010110000000000,
    17'b00010110011110110,
    17'b00010111110101110,
    17'b00011001110000101,
    17'b00011101010001111,
    17'b00011111111010111,
    17'b00100010111000011,
    17'b00100110000101001,
    17'b00100111100110011,
    17'b00101010100011111,
    17'b00101101110101110,
    17'b00110100101110001,
    17'b00110100010100100,
    17'b00110100010100100,
    17'b00111000101110001,
    17'b00111011000010100,
    17'b00110111110101110,
    17'b00110101110000101,
    17'b00110111110101110,
    17'b00110111001100110,
    17'b00110010010100100,
    17'b00110100110011010,
    17'b00110101101011100,
    17'b00110110001010010,
    17'b00110101100001010,
    17'b00110100111101100,
    17'b00110111010001111,
    17'b00101001111010111,
    17'b00100101000010100,
    17'b00011110101001000,
    17'b00011010000101001,
    17'b00100001111010111,
    17'b00100000111000011,
    17'b00011100000101001,
    17'b00011001111010111,
    17'b00100101101011100,
    17'b00111101011100001,
    17'b01001001100001010,
    17'b01000110111101100,
    17'b01000010110011010,
    17'b00111110101110001,
    17'b00111000111000011,
    17'b00110000000101001,
    17'b00101011111010111,
    17'b00101010011001101,
    17'b00101010101001000,
    17'b00101100011001101,
    17'b00110001010001111,
    17'b00110101010111000,
    17'b00111000011001101,
    17'b00111010000000000,
    17'b00111001100001010,
    17'b00111000011110110,
    17'b00110111110101110,
    17'b00110111010001111,
    17'b00110110110011010,
    17'b00111000111000011,
    17'b00110110001010010,
    17'b00110111000111101,
    17'b00111000001010010,
    17'b00101101011100001,
    17'b00101110001010010,
    17'b00101101010111000,
    17'b00101011110000101,
    17'b00101100011001101,
    17'b00101110011110110,
    17'b00101100110011010,
    17'b00101011010001111,
    17'b00100111100110011,
    17'b00100110000101001,
    17'b00100111000111101,
    17'b00101010110011010,
    17'b00101011000010100,
    17'b00101101100110011,
    17'b00111000101001000,
    17'b00111001011100001,
    17'b00111111001100110,
    17'b01000000001111011,
    17'b01000000010100100,
    17'b00111110011001101,
    17'b01000000100011111,
    17'b00111101001100110,
    17'b01000001000010100,
    17'b01000010101001000,
    17'b00111011111010111,
    17'b00111101110000101,
    17'b00111001011100001,
    17'b00110101010001111,
    17'b00110000000000000,
    17'b00101100010100100,
    17'b00101010010100100,
    17'b00101001010111000,
    17'b00100111010111000,
    17'b00100101101011100,
    17'b00100110010100100,
    17'b00100101110000101,
    17'b00100101001100110,
    17'b00101010111101100,
    17'b00100011110101110,
    17'b00011010111101100,
    17'b00011000001010010,
    17'b00010111100001010,
    17'b00011001010001111,
    17'b00011101100110011,
    17'b00011100011110110,
    17'b00100001011100001,
    17'b00100111100110011,
    17'b00101011011100001,
    17'b00110011000010100,
    17'b00110111010111000,
    17'b00111001011100001,
    17'b00111010010100100,
    17'b00111010011001101,
    17'b00111100011001101,
    17'b00111010000000000,
    17'b00110101100001010,
    17'b00110001110000101,
    17'b00110000000101001,
    17'b00110000111000011,
    17'b00110011010111000,
    17'b00111000011001101,
    17'b00111000001111011,
    17'b01000000000101001,
    17'b01001000000101001,
    17'b01001100101110001,
    17'b01001110101110001,
    17'b01001011010111000,
    17'b01000110010100100,
    17'b00111111111010111,
    17'b00111100000000000,
    17'b00111010011001101,
    17'b00110111011100001,
    17'b00110101000111101,
    17'b00110011111010111,
    17'b00110010011001101,
    17'b00101111100001010,
    17'b00101101110101110,
    17'b00101011110000101,
    17'b00101001001100110,
    17'b00100110001111011,
    17'b00100011111010111,
    17'b00100001100110011,
    17'b00011111100110011,
    17'b00011101100110011,
    17'b00011011110000101,
    17'b00011011000010100,
    17'b00011011000010100,
    17'b00011011100001010,
    17'b00011100101001000,
    17'b00011101010111000,
    17'b00011101001100110,
    17'b00011011111010111,
    17'b00011100000101001,
    17'b00011010111101100,
    17'b00100010101001000,
    17'b00011110000101001,
    17'b00011010000000000,
    17'b00100000011110110,
    17'b00100011100110011,
    17'b00100100011001101,
    17'b00100100011110110,
    17'b00100100110011010,
    17'b00100111100110011,
    17'b00101011001100110,
    17'b00101111001100110,
    17'b00110101100110011,
    17'b00111101100110011,
    17'b01010011110101110,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01111111111111111,
    17'b01101001011100001,
    17'b00110001110000101,
    17'b11111101111010111,
    17'b11100101100110011,
    17'b11001110001111011,
    17'b10101111110101110,
    17'b10110011000010100,
    17'b11100001100001010,
    17'b00010011101011100,
    17'b00110000110011010,
    17'b00111011000010100,
    17'b01000100111101100,
    17'b01011011000111101,
    17'b01010111101011100,
    17'b01001010100011111,
    17'b01000010100011111,
    17'b01000000111000011,
    17'b01000001100110011,
    17'b01000001110101110,
    17'b01000001111010111,
    17'b01000000110011010,
    17'b00111100101110001,
    17'b00111010111000011,
    17'b00111001011100001,
    17'b00111000100011111,
    17'b00110111101011100,
    17'b00110111001100110,
    17'b00111000011110110,
    17'b00111000111101100,
    17'b00111000111101100,
    17'b00111001001100110,
    17'b00111000101110001,
    17'b00111000110011010,
    17'b00110111011100001,
    17'b00110111011100001,
    17'b00110110010100100,
    17'b00110110101110001,
    17'b00110101011100001,
    17'b00110100100011111,
    17'b00110100001111011,
    17'b00110101100001010,
    17'b00110101110000101,
    17'b00110110000000000,
    17'b00110101110101110,
    17'b00110110011110110,
    17'b00111000011001101,
    17'b00110111101011100,
    17'b00111000001010010,
    17'b00111001010111000,
    17'b00111010011001101,
    17'b00111100011001101,
    17'b00111100111101100,
    17'b00111101100001010,
    17'b00111110010100100,
    17'b00111110110011010,
    17'b00111110001111011,
    17'b00111101010001111,
    17'b00111100001010010,
    17'b00111010111101100,
    17'b00111001100001010,
    17'b00111000010100100,
    17'b00110111100001010,
    17'b00110110100011111,
    17'b00110101100110011,
    17'b00110100010100100,
    17'b00110011000111101,
    17'b00110001110000101,
    17'b00110000000000000,
    17'b00101101100110011,
    17'b00101100000000000,
    17'b00101010101001000,
    17'b00101001010111000,
    17'b00100111110101110,
    17'b00100110001010010,
    17'b00100100001111011,
    17'b00100010010100100,
    17'b00100000111000011,
    17'b00100000111101100,
    17'b00100001100001010,
    17'b00100010011001101,
    17'b00100011100001010,
    17'b00100101011100001,
    17'b00100101100110011,
    17'b00100111101011100,
    17'b00101001001100110,
    17'b00101000111000011,
    17'b00101000000000000,
    17'b00100111110101110,
    17'b00101000000000000,
    17'b00100111101011100,
    17'b00100110111000011,
    17'b00100110010100100,
    17'b00100110110011010,
    17'b00100100000000000,
    17'b00100000011110110,
    17'b00011111000010100,
    17'b00011111000010100,
    17'b00011111000010100,
    17'b00100000001010010,
    17'b00011010001111011,
    17'b00011000110011010,
    17'b00011000011001101,
    17'b00011011100001010,
    17'b00011000000000000,
    17'b00010110000101001,
    17'b00010111100001010,
    17'b00010110100011111,
    17'b00100001111010111,
    17'b00100011110000101,
    17'b00010110011001101,
    17'b00001101000111101,
    17'b00010100000101001,
    17'b00011000001010010,
    17'b00010110000101001,
    17'b00010100001111011,
    17'b00010011000111101,
    17'b00010100111000011,
    17'b00010110110011010,
    17'b00011000000000000,
    17'b00011001010111000,
    17'b00011010111000011,
    17'b00011100101001000,
    17'b00011101101011100,
    17'b00011110011001101,
    17'b00011111000010100,
    17'b00011111001100110,
    17'b00011110101110001,
    17'b00011110000101001,
    17'b00011101001100110,
    17'b00011011110000101,
    17'b00011010111000011,
    17'b00011010000000000,
    17'b00011001010111000,
    17'b00011001010111000,
    17'b00011001001100110,
    17'b00011000110011010,
    17'b00011000001010010,
    17'b00010110101001000,
    17'b00010101011100001,
    17'b00010100000101001,
    17'b00010010111000011,
    17'b00010001011100001,
    17'b00010000011001101,
    17'b00001111001100110,
    17'b00001110011110110,
    17'b00001110000101001,
    17'b00001101111010111,
    17'b00001110000000000,
    17'b00001110011110110,
    17'b00001110111000011,
    17'b00001110110011010,
    17'b00001110111101100,
    17'b00001111000111101,
    17'b00001111000010100,
    17'b00001110110011010,
    17'b00001101110101110,
    17'b00001100000000000,
    17'b00001001111010111,
    17'b00001001010001111,
    17'b00001001011100001,
    17'b00001011010001111,
    17'b00001110011110110,
    17'b00010100110011010,
    17'b00100101100001010,
    17'b00100011100001010,
    17'b00011100111000011,
    17'b00011110000000000,
    17'b00011111110000101,
    17'b00100010001111011,
    17'b00100101001100110,
    17'b00100110011110110,
    17'b00100111101011100,
    17'b00101000100011111,
    17'b00101001111010111,
    17'b00101001101011100,
    17'b00101001011100001,
    17'b00101001001100110,
    17'b00101000100011111,
    17'b00100110110011010,
    17'b00100101111010111,
    17'b00100110011110110,
    17'b00100110100011111,
    17'b00100101111010111,
    17'b00100101110000101,
    17'b00100101110000101,
    17'b00100110001010010,
    17'b00100110111101100,
    17'b00101000111000011,
    17'b00101010011001101,
    17'b00101011000111101,
    17'b00101011010001111,
    17'b00101100100011111,
    17'b00110010001111011,
    17'b00110100101110001,
    17'b00110110000000000,
    17'b00110100011110110,
    17'b00101010011110110,
    17'b00110000011001101,
    17'b00110001100001010,
    17'b00110010001111011,
    17'b00110010011110110,
    17'b00110011000111101,
    17'b00110100010100100,
    17'b00110100110011010,
    17'b00110110000000000,
    17'b00110000111000011,
    17'b00110010010100100,
    17'b00110001100001010,
    17'b00110000111101100,
    17'b00101101110101110,
    17'b00101010100011111,
    17'b00100011100001010,
    17'b00011110110011010,
    17'b00011010111000011,
    17'b00010110110011010,
    17'b00010001001100110,
    17'b00001101011100001,
    17'b00001011010001111,
    17'b00001000001111011,
    17'b00000110101110001,
    17'b00000110101001000,
    17'b00000110000000000,
    17'b00000101100110011,
    17'b00000101001100110,
    17'b00000100101001000,
    17'b00000011110000101,
    17'b00000011010001111,
    17'b00000010111101100,
    17'b00000011001100110,
    17'b00000011000111101,
    17'b00000010111000011,
    17'b00000010111000011,
    17'b00000011001100110,
    17'b00000011100001010,
    17'b00000011100001010,
    17'b00000011000111101,
    17'b00000010101001000,
    17'b00000001101011100,
    17'b00000100000000000,
    17'b00000101100110011,
    17'b11111010111101100,
    17'b11111110000101001,
    17'b11111111010111000,
    17'b00000001100110011,
    17'b11111111001100110,
    17'b11111100000101001,
    17'b11111000101110001,
    17'b11110100010100100,
    17'b11110011010001111,
    17'b11101110011001101,
    17'b11101001101011100,
    17'b11100111001100110,
    17'b11100101001100110,
    17'b11100010101001000,
    17'b11100001011100001,
    17'b11011110011110110,
    17'b11011100110011010,
    17'b11011010101001000,
    17'b11011010011110110,
    17'b11011000111000011,
    17'b11011000010100100,
    17'b11010110111101100,
    17'b11001011100110011,
    17'b11001011000010100,
    17'b11001101010111000,
    17'b11001111000010100,
    17'b11001111010111000,
    17'b11001110101001000,
    17'b11001101000111101,
    17'b11001100000101001,
    17'b11001011001100110,
    17'b11001001111010111,
    17'b11001000110011010,
    17'b11000111010111000,
    17'b11000101101011100,
    17'b11000011000010100,
    17'b11000000111000011,
    17'b10111110100011111,
    17'b10111100000000000,
    17'b10111010000101001,
    17'b10111010100011111,
    17'b10111011110000101,
    17'b10111100001010010,
    17'b10111100000000000,
    17'b10111100011001101,
    17'b10111100010100100,
    17'b10110110111101100,
    17'b10101110111000011,
    17'b10100110101110001,
    17'b10100010010100100,
    17'b10100010001111011,
    17'b10100100101110001,
    17'b10100111110101110,
    17'b10101001111010111,
    17'b10101010000101001,
    17'b10101001101011100,
    17'b10101001101011100,
    17'b10101010000101001,
    17'b10101010110011010,
    17'b10101011111010111,
    17'b10101101010111000,
    17'b10101110001010010,
    17'b10100111001100110,
    17'b10100011100110011,
    17'b10100001001100110,
    17'b10011111000010100,
    17'b10011101110000101,
    17'b10011101100110011,
    17'b10011110100011111,
    17'b10100010000000000,
    17'b10100010101001000,
    17'b10100000101001000,
    17'b10011110011110110,
    17'b10011101010111000,
    17'b10011101101011100,
    17'b10011110001111011,
    17'b10011111011100001,
    17'b10100000011110110,
    17'b10100001000111101,
    17'b10100001010111000,
    17'b10100001010001111,
    17'b10100001011100001,
    17'b10100010000101001,
    17'b10100001011100001,
    17'b10100000111000011,
    17'b10100000011110110,
    17'b10011111110101110,
    17'b10011111010111000,
    17'b10011111010001111,
    17'b10011110111000011,
    17'b10011110011110110,
    17'b10011110001010010,
    17'b10011101100001010,
    17'b10011101110101110,
    17'b10011010001010010,
    17'b10011010011001101,
    17'b10011010000000000,
    17'b10011010111000011,
    17'b10011011000010100,
    17'b10011100000000000,
    17'b10011100111101100,
    17'b10010100010100100,
    17'b10000000000000000,
    17'b10000000000000000,
    17'b10000001110101110,
    17'b10001101001100110,
    17'b10011001011100001,
    17'b10100001110000101,
    17'b10011101101011100,
    17'b10011100000000000,
    17'b10011011011100001,
    17'b10011101100110011,
    17'b10100100000000000,
    17'b10101101000010100,
    17'b10100100001111011,
    17'b10100110011110110,
    17'b10100101111010111,
    17'b10100011101011100,
    17'b10100010011110110,
    17'b10100100001111011,
    17'b10100110011001101,
    17'b10101100111000011,
    17'b10110001010111000,
    17'b10110101000010100,
    17'b10111000100011111,
    17'b10111100010100100,
    17'b11000001110000101,
    17'b11001001011100001,
    17'b11101000111101100,
    17'b11101100111101100,
    17'b11101111110101110,
    17'b11110010010100100,
    17'b11110100011110110,
    17'b11110101010111000,
    17'b11110110000101001,
    17'b11110110011001101,
    17'b11110111110101110,
    17'b11111010000000000,
    17'b11111011110000101,
    17'b11111110000101001,
    17'b00000000111000011,
    17'b00000011100110011,
    17'b00000111101011100,
    17'b00001011110101110,
    17'b00010000000000000,
    17'b00010011011100001,
    17'b00010111000010100,
    17'b00011100000000000,
    17'b00011110100011111,
    17'b00100000001111011,
    17'b00100001010001111,
    17'b00100001111010111,
    17'b00100010000000000,
    17'b00100001010001111,
    17'b00100000010100100,
    17'b00011111111010111,
    17'b00011111110101110,
    17'b00100000011110110,
    17'b00100000101001000,
    17'b00100000000101001,
    17'b00100000000000000,
    17'b00011111010001111,
    17'b00011111000111101,
    17'b00100000001010010,
    17'b00100000111000011,
    17'b00100001000111101,
    17'b00100010000101001,
    17'b00100010101110001,
    17'b00100010001111011,
    17'b00100010000000000,
    17'b00100011100110011,
    17'b00100101001100110,
    17'b00100101010111000,
    17'b00100101011100001,
    17'b00101001110101110,
    17'b00101011110101110,
    17'b00101110101001000,
    17'b00110010101110001,
    17'b00110110010100100,
    17'b00111100101110001,
    17'b00111011100110011,
    17'b00111111001100110,
    17'b01000100101110001,
    17'b01000110001111011,
    17'b01001000100011111,
    17'b01001101010001111,
    17'b01001110000101001,
    17'b01001111101011100,
    17'b01010011100110011,
    17'b01010000100011111,
    17'b01001110011110110,
    17'b01001100111000011,
    17'b01001000110011010,
    17'b01000101100001010,
    17'b01000011000111101,
    17'b00111111011100001,
    17'b00111011010001111,
    17'b00110111001100110,
    17'b00110010110011010,
    17'b00101111100001010,
    17'b00101011011100001,
    17'b00100100111000011,
    17'b00100011000010100,
    17'b00100010011001101,
    17'b00100001000010100,
    17'b00011110111000011,
    17'b00011111100110011,
    17'b00100001000010100,
    17'b00100000100011111,
    17'b00011111000010100,
    17'b00011101111010111,
    17'b00011101111010111,
    17'b00011011101011100,
    17'b00011101101011100,
    17'b00100011000010100,
    17'b00100111011100001,
    17'b00100100011001101,
    17'b00011111110101110,
    17'b00011110000000000,
    17'b00011100111000011,
    17'b00011010000000000,
    17'b00010111010111000,
    17'b00010100001010010,
    17'b00010000001111011,
    17'b00001011000010100,
    17'b00000111110101110,
    17'b00000101001100110,
    17'b00000010001111011,
    17'b11111110010100100,
    17'b11111100010100100,
    17'b11111010001111011,
    17'b11111000100011111,
    17'b11110101111010111,
    17'b11110100001111011,
    17'b11110011110101110,
    17'b11110011110101110,
    17'b11110000101001000,
    17'b11101110100011111,
    17'b11101110110011010,
    17'b11101010101110001,
    17'b11100111100110011,
    17'b11101101110101110,
    17'b11101100110011010,
    17'b11011100010100100,
    17'b11011010100011111,
    17'b11001111010001111,
    17'b11010111011100001,
    17'b11100110001111011,
    17'b11101111000111101,
    17'b11101100100011111,
    17'b11101011000010100,
    17'b11101001010001111,
    17'b11100111011100001,
    17'b11100010011001101,
    17'b11100000010100100,
    17'b11100000101110001,
    17'b11011110101001000,
    17'b11011011101011100,
    17'b11011000110011010,
    17'b11010110101110001,
    17'b11010100111101100,
    17'b11010011000111101,
    17'b11010000111000011,
    17'b11001111000111101,
    17'b11001110000000000,
    17'b11001101100110011,
    17'b11001110011001101,
    17'b11001110011110110,
    17'b11001110001010010,
    17'b11001110001010010,
    17'b11001100111000011,
    17'b11001010010100100,
    17'b11000111001100110,
    17'b11000011010001111,
    17'b11000000010100100,
    17'b10111110111101100,
    17'b10111111110000101,
    17'b10111110110011010,
    17'b10111011110000101,
    17'b10111000011001101,
    17'b10110110111101100,
    17'b10110110010100100,
    17'b10110110010100100,
    17'b10110111101011100,
    17'b10111001000111101,
    17'b10111001000010100,
    17'b10111001010111000,
    17'b10111010010100100,
    17'b10111011010001111,
    17'b10111010101001000,
    17'b10111001100001010,
    17'b10111000101001000,
    17'b10110111110101110,
    17'b10110111100001010,
    17'b10110110101110001,
    17'b10110111000010100,
    17'b10110110011110110,
    17'b10110110000000000,
    17'b10110101011100001,
    17'b10110101101011100,
    17'b10110101100001010,
    17'b10110101110000101,
    17'b10110100110011010,
    17'b10110011110000101,
    17'b10110010011110110,
    17'b10110010000101001,
    17'b10110001110000101,
    17'b10110001100001010,
    17'b10110001110101110,
    17'b10110011100001010,
    17'b10110111000111101,
    17'b10110111010001111,
    17'b10110100000101001,
    17'b10111010001010010,
    17'b10111001111010111,
    17'b10111101000010100,
    17'b10110100101110001,
    17'b10110001010001111,
    17'b10111000111101100,
    17'b10110010111000011,
    17'b10110011110000101,
    17'b10110101110101110,
    17'b10101111110000101,
    17'b10110100000000000,
    17'b10110010001111011,
    17'b10110110011001101,
    17'b10101011110000101,
    17'b10101101111010111,
    17'b10110001100110011,
    17'b10111111001100110,
    17'b10111010101110001,
    17'b10111000101110001,
    17'b10111001110101110,
    17'b10111000011001101,
    17'b10110101111010111,
    17'b10110110000101001,
    17'b10111001000010100,
    17'b10110110011001101,
    17'b10110100011001101,
    17'b10110011100001010,
    17'b10110011100001010,
    17'b10110001010001111,
    17'b10110001101011100,
    17'b10110010011001101,
    17'b10110110000101001,
    17'b10110111100110011,
    17'b10111001000010100,
    17'b10111001110000101,
    17'b10111011001100110,
    17'b10111100101110001,
    17'b10111101110000101,
    17'b10111110110011010,
    17'b11000000100011111,
    17'b11000010100011111,
    17'b11000010110011010,
    17'b11000011110101110,
    17'b11000111010001111,
    17'b11001001110101110,
    17'b11001100011001101,
    17'b11001111101011100,
    17'b11010001000010100,
    17'b11010001100110011,
    17'b11010001110101110,
    17'b11010010111101100,
    17'b11010100101110001,
    17'b11010101000010100,
    17'b11010110000000000,
    17'b11011000010100100,
    17'b11011001110101110,
    17'b11011010101110001,
    17'b11011011000111101,
    17'b11011001111010111,
    17'b11011010010100100,
    17'b11011011111010111,
    17'b11011110010100100,
    17'b11100001110101110,
    17'b11100101000010100,
    17'b11100110001111011,
    17'b11100111001100110,
    17'b11100111110000101,
    17'b11100111111010111,
    17'b11101000000101001,
    17'b11101000001111011,
    17'b11101001000111101,
    17'b11101010100011111,
    17'b11101101000111101,
    17'b11110000000101001,
    17'b11110001011100001,
    17'b11110010101001000,
    17'b11110101100001010,
    17'b11111010011110110,
    17'b11111101110101110,
    17'b00000000000000000,
    17'b00000001100110011,
    17'b00000100001010010,
    17'b00000110101001000,
    17'b00001000000000000,
    17'b00000111110101110,
    17'b00000111110000101,
    17'b00001000001111011,
    17'b00001000000000000,
    17'b00000111110000101,
    17'b00000111100001010,
    17'b00000110011110110,
    17'b00000110000000000,
    17'b00000110101001000,
    17'b00000111010001111,
    17'b00000111101011100,
    17'b00000110101110001,
    17'b00000101010001111,
    17'b00000100001010010,
    17'b00000010110011010,
    17'b00000000111000011,
    17'b00000000001010010,
    17'b00000000111000011,
    17'b00000010100011111,
    17'b00000100101110001,
    17'b00010111000010100,
    17'b00011100101110001,
    17'b00011111100001010,
    17'b00100101111010111,
    17'b00101100100011111,
    17'b00110001010111000,
    17'b00110100011001101,
    17'b00111000011001101,
    17'b00111100000000000,
    17'b00111101010001111,
    17'b00111101101011100,
    17'b00111110010100100,
    17'b00111111110000101,
    17'b00111111110000101,
    17'b00111111101011100,
    17'b00111111101011100,
    17'b01000000000000000,
    17'b01000000001111011,
    17'b01000000011001101,
    17'b01000000001111011,
    17'b01000000000000000,
    17'b01000000011110110,
    17'b00111111011100001,
    17'b00111101110101110,
    17'b00111100101001000,
    17'b00111010111000011,
    17'b00111000101110001,
    17'b00110111001100110,
    17'b00110101100001010,
    17'b00110100000101001,
    17'b00110001100110011,
    17'b00110000111000011,
    17'b00101111100110011,
    17'b00101100100011111,
    17'b00101010101001000,
    17'b00101010000101001,
    17'b00101000110011010,
    17'b00100110111101100,
    17'b00100101101011100,
    17'b00100100110011010,
    17'b00100011111010111,
    17'b00100011010111000,
    17'b00100010011110110,
    17'b00100010011001101,
    17'b00100010001111011,
    17'b00100010000101001,
    17'b00100001101011100,
    17'b00100001011100001,
    17'b00100010011001101,
    17'b00100010110011010,
    17'b00100010111101100,
    17'b00100011100001010,
    17'b00100011110000101,
    17'b00100011011100001,
    17'b00100011011100001,
    17'b00100011111010111,
    17'b00100001110000101,
    17'b00100000011001101,
    17'b00100000000101001,
    17'b00010110110011010,
    17'b00010101000010100,
    17'b00010010000101001,
    17'b00010000101001000,
    17'b00001111100110011,
    17'b00001111000010100,
    17'b00001110111101100,
    17'b00001110101110001,
    17'b00001101001100110,
    17'b00001100001111011,
    17'b00001011000111101,
    17'b00001001100110011,
    17'b00001000001010010,
    17'b00000110011001101,
    17'b00000101111010111,
    17'b00000010111101100,
    17'b00000000010100100,
    17'b11111110101001000,
    17'b11111100101110001,
    17'b11111011001100110,
    17'b11111010011001101,
    17'b11111001010111000,
    17'b11111001001100110,
    17'b11111001100001010,
    17'b11111010011110110,
    17'b11111010111101100,
    17'b11111011010001111,
    17'b11111011010001111,
    17'b11111010001010010,
    17'b11111000111101100,
    17'b11110111110101110,
    17'b11110110011110110,
    17'b11110100101110001,
    17'b11110011000111101,
    17'b11110000110011010,
    17'b11101110011001101,
    17'b11101011001100110,
    17'b11101000111000011,
    17'b11100110101001000,
    17'b11100100011110110,
    17'b11100001001100110,
    17'b11011111000010100,
    17'b11011101100001010,
    17'b11011011111010111,
    17'b11011010110011010,
    17'b11011010010100100,
    17'b11011010011001101,
    17'b11011010101110001,
    17'b11011111101011100,
    17'b11100000101110001,
    17'b11100010011110110,
    17'b11100111011100001,
    17'b11101100011110110,
    17'b11101001110000101,
    17'b11101110001111011,
    17'b11110010011001101,
    17'b11111001101011100,
    17'b00100001010001111,
    17'b00011101001100110,
    17'b10000000000000000,
    17'b10001111010111000,
    17'b10100110001111011,
    17'b10101100011110110,
    17'b11000010111101100,
    17'b11001000111000011,
    17'b11001010111101100,
    17'b11001101001100110,
    17'b11001011001100110,
    17'b11001001011100001,
    17'b11001010101001000,
    17'b11001101010001111,
    17'b11001110011001101,
    17'b11001111100110011,
    17'b11001111000010100,
    17'b11001100001010010,
    17'b11001001110000101,
    17'b11000111100001010,
    17'b11000101010001111,
    17'b11000011010001111,
    17'b11000010000000000,
    17'b11000001000111101,
    17'b11000001000010100,
    17'b11000010000000000,
    17'b11000010011110110,
    17'b11000011010001111,
    17'b11000100000000000,
    17'b11001000100011111,
    17'b11001001011100001,
    17'b11001010001010010,
    17'b11001011000010100,
    17'b11001011101011100,
    17'b11001011101011100,
    17'b11001011101011100,
    17'b11001011011100001,
    17'b11001010111000011,
    17'b11001010010100100,
    17'b11001010000000000,
    17'b11001001101011100,
    17'b11001010000101001,
    17'b11001010101001000,
    17'b11001010110011010,
    17'b11001010111000011,
    17'b11001010101001000,
    17'b11001001001100110,
    17'b11000111101011100,
    17'b11000101100001010,
    17'b11000011110101110,
    17'b11000011001100110,
    17'b11000010110011010,
    17'b11000010001111011,
    17'b11000010100011111,
    17'b11000010111101100,
    17'b11000011001100110,
    17'b11000011010111000,
    17'b11000011000111101,
    17'b11000010101110001,
    17'b11000010001111011,
    17'b11000010000000000,
    17'b11000010000000000,
    17'b11000010000101001,
    17'b11000010111000011,
    17'b11000011010111000,
    17'b11000100001111011,
    17'b11000100101110001,
    17'b11000101111010111,
    17'b11001101110000101,
    17'b11010001001100110,
    17'b11010110001010010,
    17'b11011011101011100,
    17'b11100001110000101,
    17'b11101000111101100,
    17'b11110000101110001,
    17'b11110110011001101,
    17'b11111100000000000,
    17'b00000011001100110,
    17'b00000111101011100,
    17'b00001011100001010,
    17'b00001111001100110,
    17'b00010011110101110,
    17'b00010110101001000,
    17'b00011000011110110,
    17'b00011010101001000,
    17'b00011100011110110,
    17'b00011110011110110,
    17'b00011111100001010,
    17'b00100000110011010,
    17'b00100010111000011,
    17'b00100100101001000,
    17'b00100110111101100,
    17'b00101001100110011,
    17'b00101011100110011,
    17'b00101101100001010,
    17'b00101111011100001,
    17'b00101111011100001,
    17'b00101110001010010,
    17'b00101101001100110,
    17'b00101100111000011,
    17'b00101110000000000,
    17'b00101110111101100,
    17'b00110000000101001,
    17'b00110000010100100,
    17'b00101111100001010,
    17'b00101111101011100,
    17'b00110000001111011,
    17'b00110000011001101,
    17'b00110000010100100,
    17'b00110000101001000,
    17'b00110000011001101,
    17'b00101111100001010,
    17'b00101111100110011,
    17'b00101110010100100,
    17'b00101110101001000,
    17'b00101110001111011,
    17'b00101111010001111,
    17'b00101110001010010,
    17'b00101111100001010,
    17'b00101111011100001,
    17'b00110000101001000,
    17'b00110010011110110,
    17'b00110011100001010,
    17'b00110101011100001,
    17'b00110100111101100,
    17'b00110101110000101,
    17'b00110100001111011,
    17'b00110101100110011,
    17'b00110110101001000,
    17'b00110110111000011,
    17'b00110111011100001,
    17'b00110111000111101,
    17'b00110110111101100,
    17'b00110111011100001,
    17'b00110111010001111,
    17'b00110110111101100,
    17'b00110110000000000,
    17'b00110101010001111,
    17'b00110111000111101,
    17'b00111000111000011,
    17'b00111010001010010,
    17'b00111100001010010,
    17'b00111011011100001,
    17'b00111001100110011,
    17'b00110111101011100,
    17'b00111011000010100,
    17'b00111100101001000,
    17'b00111110000000000,
    17'b00111100011001101,
    17'b00111111010111000,
    17'b00111111110000101,
    17'b01000000011110110,
    17'b01000000100011111,
    17'b00111111111010111,
    17'b00111110111000011,
    17'b00111110111000011,
    17'b00111110011001101,
    17'b00111110011110110,
    17'b00111110101110001,
    17'b00111100111101100,
    17'b00111011110101110,
    17'b00110001100001010,
    17'b00011101010001111,
    17'b00010100110011010,
    17'b00110000111101100,
    17'b00011010101110001,
    17'b00011010001111011,
    17'b00100101010001111,
    17'b00110011110101110,
    17'b01000010111000011,
    17'b01001011101011100,
    17'b01001010110011010,
    17'b01001101101011100,
    17'b01010001000111101,
    17'b01010000001111011,
    17'b01001110100011111,
    17'b01001101110101110,
    17'b01001100010100100,
    17'b01001010110011010,
    17'b01001000011110110,
    17'b01000100110011010,
    17'b00111111011100001,
    17'b00111100100011111,
    17'b00111010011001101,
    17'b00111000011110110,
    17'b00110110111000011,
    17'b00110101011100001,
    17'b00110100011110110,
    17'b00110011001100110,
    17'b00110010101110001,
    17'b00110001110101110,
    17'b00101101110101110,
    17'b00101011101011100,
    17'b00101100101110001,
    17'b00101110011001101,
    17'b00110000101001000,
    17'b00110010011110110,
    17'b00110100000101001,
    17'b00110101000010100,
    17'b00110110000000000,
    17'b00110110010100100,
    17'b00110110010100100,
    17'b00110110000000000,
    17'b00110101000010100,
    17'b00110100000101001,
    17'b00110100011110110,
    17'b00110100111000011,
    17'b00110101000010100,
    17'b00110101011100001,
    17'b00110110010100100,
    17'b00110110110011010,
    17'b00110111100001010,
    17'b00111000001010010,
    17'b00111001010111000,
    17'b00111010011110110,
    17'b01001010000101001,
    17'b01010100111000011,
    17'b01000001100110011,
    17'b00110110010100100,
    17'b00110011100001010,
    17'b00110000000101001,
    17'b00101100010100100,
    17'b00101001111010111,
    17'b00101000100011111,
    17'b00100111100001010,
    17'b00100110001010010,
    17'b00100110000000000,
    17'b00100110001010010,
    17'b00100110111000011,
    17'b00100111111010111,
    17'b00101001010111000,
    17'b00101010000000000,
    17'b00101010100011111,
    17'b00101011100110011,
    17'b00101100011001101,
    17'b00101100101110001,
    17'b00101100101001000,
    17'b00101100111000011,
    17'b00101101100001010,
    17'b00101101101011100,
    17'b00101101110000101,
    17'b00101101100110011,
    17'b00101101011100001,
    17'b00101100110011010,
    17'b00101011110000101,
    17'b00101010101110001,
    17'b00101001110000101,
    17'b00101010110011010,
    17'b00101010110011010,
    17'b00101010101110001,
    17'b00101011000010100,
    17'b00101011111010111,
    17'b00101100010100100,
    17'b00101100110011010,
    17'b00101101001100110,
    17'b00101100111000011,
    17'b00101100111000011,
    17'b00101101010001111,
    17'b00101101100110011,
    17'b00101101110000101,
    17'b00101101100001010,
    17'b00101101011100001,
    17'b00101101001100110,
    17'b00101101000010100,
    17'b00101101111010111,
    17'b00101110110011010,
    17'b00101111001100110,
    17'b00101111011100001,
    17'b00101111010111000,
    17'b00101111000010100,
    17'b00101110111000011,
    17'b00101110101110001,
    17'b00101110000000000,
    17'b00101101000010100,
    17'b00101100000101001,
    17'b00101011100110011,
    17'b00101010111101100,
    17'b00101010010100100,
    17'b00101001110101110,
    17'b00101001101011100,
    17'b00101001100001010,
    17'b00101001100110011,
    17'b00101001111010111,
    17'b00101010000101001,
    17'b00101010000000000,
    17'b00101001000010100,
    17'b00100111110000101,
    17'b00100110100011111,
    17'b00100101110000101,
    17'b00100101001100110,
    17'b00100100111101100,
    17'b00100100000101001,
    17'b00100010111000011,
    17'b00100001100110011,
    17'b00100000111000011,
    17'b00100000001111011,
    17'b00011100001010010,
    17'b00011011100110011,
    17'b00011011000111101,
    17'b00011010101110001,
    17'b00011010000101001,
    17'b00011001011100001,
    17'b00011000101110001,
    17'b00011000000101001,
    17'b00010111000111101,
    17'b00010110101110001,
    17'b00010110101001000,
    17'b00010110101110001,
    17'b00010110101110001,
    17'b00010110101110001,
    17'b00010110101110001,
    17'b00010110111101100,
    17'b00010111001100110,
    17'b00010110111101100,
    17'b00010110101110001,
    17'b00010110000101001,
    17'b00010101100110011,
    17'b00010101000111101,
    17'b00010100100011111,
    17'b00010011011100001,
    17'b00010010100011111,
    17'b00010001100001010,
    17'b00010000011001101,
    17'b00001111000111101,
    17'b00001110001111011,
    17'b00001101010111000,
    17'b00001100100011111,
    17'b00001011010111000,
    17'b00001010100011111,
    17'b00001010000101001,
    17'b00001001111010111,
    17'b00001001100110011,
    17'b00001000111101100,
    17'b00000101110000101,
    17'b00000011101011100,
    17'b00000110111000011,
    17'b00001001000010100,
    17'b00001001010111000,
    17'b00000101100001010,
    17'b00000100111101100,
    17'b00000011111010111,
    17'b00000010101001000,
    17'b00000001100110011,
    17'b00000000111000011,
    17'b00000000011001101,
    17'b11111110111101100,
    17'b11111101110101110,
    17'b11111110000000000,
    17'b11111101111010111,
    17'b11111101001100110,
    17'b11111101000010100,
    17'b11111100101110001,
    17'b11111011111010111,
    17'b11111010110011010,
    17'b11111010011110110,
    17'b11111010000000000,
    17'b11111001000111101,
    17'b11111000011001101,
    17'b11110111100110011,
    17'b11110110011110110,
    17'b11110101100110011,
    17'b11110101000010100,
    17'b11110100011110110,
    17'b11110100001010010,
    17'b11110011110000101,
    17'b11110011010111000,
    17'b11110010111101100,
    17'b11110010110011010,
    17'b11110010000000000,
    17'b11110001010001111,
    17'b11110000111000011,
    17'b11110000001010010,
    17'b11101111110101110,
    17'b11101111010001111,
    17'b11101110001010010,
    17'b11101101010111000,
    17'b11101100111000011,
    17'b11101100010100100,
    17'b11101011001100110,
    17'b11101001100001010,
    17'b11101000010100100,
    17'b11100111100110011,
    17'b11100111110000101,
    17'b11100111100001010,
    17'b11100110101110001,
    17'b11100110001111011,
    17'b11100101110000101,
    17'b11100101000111101,
    17'b11100100111000011,
    17'b11100100001111011,
    17'b11100100000000000,
    17'b11100011100001010,
    17'b11100011001100110,
    17'b11100010111101100,
    17'b11100001110101110,
    17'b11100001000010100,
    17'b11100000011001101,
    17'b11011111110101110,
    17'b11011111000010100,
    17'b11011101111010111,
    17'b11011100011001101,
    17'b11011011110000101,
    17'b11011100000101001,
    17'b11011100001010010,
    17'b11011100110011010,
    17'b11011101010001111,
    17'b11011101100110011,
    17'b11011101100001010,
    17'b11011101011100001,
    17'b11011101011100001,
    17'b11011101000111101,
    17'b11011100111101100,
    17'b11011100100011111,
    17'b11011100000101001,
    17'b11011011101011100,
    17'b11011011000111101,
    17'b11011010110011010,
    17'b11011010000000000,
    17'b11011001011100001,
    17'b11011001000010100,
    17'b11011000100011111,
    17'b11010111110101110,
    17'b11010111100110011,
    17'b11010111000111101,
    17'b11010110111101100,
    17'b11010110111000011,
    17'b11010110101110001,
    17'b11010110011110110,
    17'b11010101100110011,
    17'b11010100101001000,
    17'b11010011111010111,
    17'b11010011010111000,
    17'b11010010011110110,
    17'b11001101100001010,
    17'b11001110101001000,
    17'b11001110011110110,
    17'b11001110101110001,
    17'b11001110111101100,
    17'b11001111001100110,
    17'b11001110111101100,
    17'b11001110011110110,
    17'b11001110101110001,
    17'b11001110110011010,
    17'b11001110101001000,
    17'b11001110101110001,
    17'b11001110010100100,
    17'b11001110001111011,
    17'b11001110000000000,
    17'b11001101100001010,
    17'b11001101100110011,
    17'b11001101010001111,
    17'b11001100111000011,
    17'b11001100101110001,
    17'b11001100101001000,
    17'b11001100111000011,
    17'b11001101001100110,
    17'b11001101010001111,
    17'b11001101110101110,
    17'b11001110101001000,
    17'b11001111010111000,
    17'b11001111100001010,
    17'b11001110111101100,
    17'b11001110010100100,
    17'b11001101000111101,
    17'b11001010101001000,
    17'b11001010100011111,
    17'b11001010011001101,
    17'b11001010001111011,
    17'b11001010001111011,
    17'b11001010000101001,
    17'b11001001101011100,
    17'b11001001001100110,
    17'b11001000101110001,
    17'b11001000011001101,
    17'b11001000101001000,
    17'b11001001001100110,
    17'b11001001011100001,
    17'b11001001101011100,
    17'b11001010000101001,
    17'b11001010000101001,
    17'b11001001110000101,
    17'b11001001010001111,
    17'b11001001000010100,
    17'b11001000111000011,
    17'b11001001000010100,
    17'b11001001010111000,
    17'b11001001110101110,
    17'b11001010101110001,
    17'b11001100001010010,
    17'b11001101010001111,
    17'b11001110010100100,
    17'b11001110111101100,
    17'b11001111110000101,
    17'b11010000000000000,
    17'b11001111110101110,
    17'b11001111010111000,
    17'b11001111000010100,
    17'b11001110101110001,
    17'b11001110001111011,
    17'b11001101101011100,
    17'b11001101001100110,
    17'b11001011111010111,
    17'b11001001100110011,
    17'b11001000100011111,
    17'b11001000011110110,
    17'b11001000100011111,
    17'b11001000001111011,
    17'b11000111011100001,
    17'b11000110001111011,
    17'b11000100110011010,
    17'b11000100010100100,
    17'b11000011101011100,
    17'b11000011110000101,
    17'b11000011101011100,
    17'b11000011011100001,
    17'b11000011001100110,
    17'b11000011100110011,
    17'b11000011110101110,
    17'b11000100000101001,
    17'b11000100001111011,
    17'b11000100010100100,
    17'b11000100001010010,
    17'b11000100010100100,
    17'b11000100000101001,
    17'b11000100000000000,
    17'b11000100101110001,
    17'b11000110000101001,
    17'b11000101100110011,
    17'b11000101000111101,
    17'b11000100101110001,
    17'b11000100001010010,
    17'b11000011110101110,
    17'b11000011100001010,
    17'b11000011010001111,
    17'b11000011000111101,
    17'b11000010011001101,
    17'b11000010000101001,
    17'b11000001110000101,
    17'b11000000101001000,
    17'b10111111101011100,
    17'b10111110101110001,
    17'b10111101000010100,
    17'b10111011001100110,
    17'b10111010011001101,
    17'b10111000011110110,
    17'b10110111000111101,
    17'b10110111000010100,
    17'b10110110111101100,
    17'b10110110101001000,
    17'b10110110101001000,
    17'b10110110011110110,
    17'b10110110001010010,
    17'b10110101010111000,
    17'b10110100001111011,
    17'b10110010100011111,
    17'b10110011110101110,
    17'b10110101110000101,
    17'b10111000011110110,
    17'b10111011010001111,
    17'b10111100011110110,
    17'b10111100110011010,
    17'b10111100010100100,
    17'b10111011110000101,
    17'b10111010011110110,
    17'b10111001101011100,
    17'b10111000010100100,
    17'b10110111010001111,
    17'b10110100011001101,
    17'b10110010000000000,
    17'b10101111101011100,
    17'b10110001011100001,
    17'b10101101010001111,
    17'b10101111100001010,
    17'b10101111010001111,
    17'b10101110011110110,
    17'b10101110001111011,
    17'b10101001010001111,
    17'b10101000000101001,
    17'b10101000000101001,
    17'b10101000001010010,
    17'b10100111100110011,
    17'b10100100000000000,
    17'b10100000111101100,
    17'b10011111010001111,
    17'b10100010000000000,
    17'b10100001110101110,
    17'b10100011000111101,
    17'b10100100001111011,
    17'b10100100111000011,
    17'b10100110111101100,
    17'b10101000100011111,
    17'b10100110001010010,
    17'b10100101011100001,
    17'b10101001000111101,
    17'b10101011100001010,
    17'b10101010101110001,
    17'b10101100011110110,
    17'b10101001001100110,
    17'b10101001000010100,
    17'b10101000011001101,
    17'b10100111111010111,
    17'b10100110010100100,
    17'b10100010111101100,
    17'b10100000000101001,
    17'b10011111100110011,
    17'b10100000101110001,
    17'b10100000101001000,
    17'b10100010010100100,
    17'b10100010000000000,
    17'b10100000101110001,
    17'b10100000101110001,
    17'b10011110110011010,
    17'b10100000001010010,
    17'b10100101000111101,
    17'b10101100000101001,
    17'b10101101000111101,
    17'b10101011010111000,
    17'b10101011110101110,
    17'b10100100000000000,
    17'b10011110000000000,
    17'b10100001010111000,
    17'b10100101110101110,
    17'b10100010001111011,
    17'b10100000001010010,
    17'b10011110001111011,
    17'b10011110110011010,
    17'b10011000110011010,
    17'b10011110010100100,
    17'b10011111000111101,
    17'b10011001110101110,
    17'b10010111011100001,
    17'b10010111100001010,
    17'b10010100010100100,
    17'b10011011010001111,
    17'b10010100111101100,
    17'b10011000110011010,
    17'b10010111000111101,
    17'b10011001101011100,
    17'b10011100111000011,
    17'b10011101100110011,
    17'b10100001000010100,
    17'b10011000110011010,
    17'b10011010011001101,
    17'b10011011111010111,
    17'b10011110001111011,
    17'b10011110000101001,
    17'b10011101101011100,
    17'b10011110000000000,
    17'b10011110000000000,
    17'b10011110000000000,
    17'b10011111000010100,
    17'b10011111000111101,
    17'b10011111010001111,
    17'b10011111101011100,
    17'b10011111111010111,
    17'b10100000011110110,
    17'b10100000101110001,
    17'b10100000001010010,
    17'b10011111000010100,
    17'b10011101100001010,
    17'b10011011001100110,
    17'b10011001001100110,
    17'b10010111000111101,
    17'b10010101100001010,
    17'b10010100010100100,
    17'b10010100101110001,
    17'b10010101010001111,
    17'b10010101100110011,
    17'b10010110110011010,
    17'b10010111110101110,
    17'b10011000110011010,
    17'b10011010011001101,
    17'b10011100001010010,
    17'b10011101011100001,
    17'b10011110111101100,
    17'b10011111100110011,
    17'b10100000000101001,
    17'b10011111100001010,
    17'b10011111000010100,
    17'b10011110101001000,
    17'b10011110001111011,
    17'b10011011111010111,
    17'b10011011100110011,
    17'b10011011000010100,
    17'b10011001011100001,
    17'b10010100110011010,
    17'b10010001110101110,
    17'b10010001110101110,
    17'b10010010101001000,
    17'b10010100000101001,
    17'b10010100101110001,
    17'b10010101000111101,
    17'b10010011000111101,
    17'b10010010010100100,
    17'b10010010001111011,
    17'b10010010101001000,
    17'b10010011110000101,
    17'b10010101110101110,
    17'b10010111100110011,
    17'b10011000101110001,
    17'b10011001010001111,
    17'b10011010000000000,
    17'b10011010010100100,
    17'b10011010110011010,
    17'b10011011011100001,
    17'b10011100000101001,
    17'b10011100101110001,
    17'b10011100111000011,
    17'b10011110001010010,
    17'b10011110111101100,
    17'b10011111001100110,
    17'b10011110111101100,
    17'b10011110001010010,
    17'b10011101011100001,
    17'b10011100101110001,
    17'b10011100000000000,
    17'b10011011100001010,
    17'b10011011011100001,
    17'b10011010101001000,
    17'b10011001000010100,
    17'b10010111010111000,
    17'b10010111101011100,
    17'b10011001001100110,
    17'b10011011000010100,
    17'b10011101110000101,
    17'b10011110111000011,
    17'b10011111001100110,
    17'b10011111000111101,
    17'b10011110111101100,
    17'b10011110101001000,
    17'b10011110111101100,
    17'b10011111010111000,
    17'b10011111110101110,
    17'b10100000001111011,
    17'b10100000101110001,
    17'b10100001000010100,
    17'b10100001011100001,
    17'b10100001110101110,
    17'b10100001111010111,
    17'b10100001110101110,
    17'b10100010000101001,
    17'b10100010001010010,
    17'b10100001111010111,
    17'b10100001101011100,
    17'b10100001111010111,
    17'b10100010011110110,
    17'b10100011001100110,
    17'b10100100001111011,
    17'b10100101000111101,
    17'b10100110001010010,
    17'b10100110110011010,
    17'b10100111010001111,
    17'b10101000001010010,
    17'b10101001100110011,
    17'b10101011000010100,
    17'b10101011011100001,
    17'b10101010111101100,
    17'b10101110000101001,
    17'b10110000100011111,
    17'b10110010101001000,
    17'b10110101000111101,
    17'b10110110000000000,
    17'b10110110110011010,
    17'b10110111110000101,
    17'b10111001001100110,
    17'b10111010011001101,
    17'b10111011100001010,
    17'b10111100110011010,
    17'b10111110101001000,
    17'b11000000011110110,
    17'b11000010000000000,
    17'b11000011100001010,
    17'b11000100001010010,
    17'b11000100110011010,
    17'b11000101100001010,
    17'b11000111000111101,
    17'b11001000101110001,
    17'b11001010101110001,
    17'b11001100101001000,
    17'b11001111000111101,
    17'b11010000111000011,
    17'b11010010010100100,
    17'b11010011100001010,
    17'b11010101000111101,
    17'b11010101111010111,
    17'b11010110011001101,
    17'b11010110101001000,
    17'b11010110101110001,
    17'b11010110101110001,
    17'b11010110001010010,
    17'b11010101110000101,
    17'b11010101100110011,
    17'b11010110001010010,
    17'b11010110111000011,
    17'b11011000001010010,
    17'b11011001010001111,
    17'b11011010011001101,
    17'b11011011101011100,
    17'b11011101010001111,
    17'b11100100000101001,
    17'b11100101110101110,
    17'b11101000000101001,
    17'b11101001110101110,
    17'b11101011110000101,
    17'b11101101100110011,
    17'b11110000000000000,
    17'b11110010000101001,
    17'b11110011110000101,
    17'b11110101100001010,
    17'b11110111111010111,
    17'b11111010000000000,
    17'b11111011101011100,
    17'b11111101010111000,
    17'b11111111000111101,
    17'b00000000000000000,
    17'b00000000111000011,
    17'b00000001100110011,
    17'b00000010101110001,
    17'b00000100000000000,
    17'b00000101000111101,
    17'b00000110011110110,
    17'b00001000001111011,
    17'b00001001001100110,
    17'b00001010001111011,
    17'b00001010111101100,
    17'b00001100001010010,
    17'b00001101100110011,
    17'b00001111000010100,
    17'b00010000100011111,
    17'b00010010000000000,
    17'b00010011001100110,
    17'b00010100000101001,
    17'b00010100111000011,
    17'b00010110101110001,
    17'b00010111110101110,
    17'b00011000101001000,
    17'b00011001110000101,
    17'b00011011000010100,
    17'b00011011111010111,
    17'b00011100111000011,
    17'b00011101011100001,
    17'b00011101110000101,
    17'b00011110011001101,
    17'b00011110110011010,
    17'b00011111010001111,
    17'b00011111100001010,
    17'b00100000010100100,
    17'b00100000111101100,
    17'b00100001110000101,
    17'b00100010000101001,
    17'b00100001101011100,
    17'b00100010001111011,
    17'b00100011000111101,
    17'b00100011100001010,
    17'b00100010101110001,
    17'b00100101100001010,
    17'b00100110001111011,
    17'b00100111010001111,
    17'b00101000011001101,
    17'b00101001110101110,
    17'b00101011000111101,
    17'b00101011010111000,
    17'b00101100001010010,
    17'b00101101000010100,
    17'b00101101100110011,
    17'b00101110000101001,
    17'b00101110011001101,
    17'b00101110001111011,
    17'b00101110000101001,
    17'b00101101101011100,
    17'b00101101000111101,
    17'b00101100001010010,
    17'b00101011101011100,
    17'b00101011110101110,
    17'b00101100011001101,
    17'b00101001100001010,
    17'b00100110101110001,
    17'b00100110000000000,
    17'b00100101111010111,
    17'b00100101010111000,
    17'b00100101001100110,
    17'b00100101000010100,
    17'b00100100111000011,
    17'b00100100100011111,
    17'b00100011110101110,
    17'b00100011001100110,
    17'b00100010011110110,
    17'b00100001111010111,
    17'b00100001110101110,
    17'b00100010011110110,
    17'b00100011110101110,
    17'b00100100101001000,
    17'b00100110000000000,
    17'b00100111100110011,
    17'b00101001100110011,
    17'b00101011100001010,
    17'b00101100111101100,
    17'b00101110000000000,
    17'b00101110010100100,
    17'b00101110010100100,
    17'b00101110101001000,
    17'b00101100111000011,
    17'b00101011000010100,
    17'b00101000111000011,
    17'b00100101111010111,
    17'b00100001001100110,
    17'b00011101110000101,
    17'b00011010011110110,
    17'b00010111010111000,
    17'b00010100011001101,
    17'b00001111110101110,
    17'b00001100010100100,
    17'b00001011100110011,
    17'b00001011110101110,
    17'b00001011100001010,
    17'b00001010110011010,
    17'b00001001001100110,
    17'b00001000010100100,
    17'b00000111001100110,
    17'b00000101100001010,
    17'b00000101110000101,
    17'b00000010011110110,
    17'b00000000000000000,
    17'b11111111000111101,
    17'b11111111110101110,
    17'b00000000110011010,
    17'b00000001000111101,
    17'b00000000010100100,
    17'b00000000101001000,
    17'b00000001001100110,
    17'b00000001110000101,
    17'b00000010100011111,
    17'b00000010100011111,
    17'b00000000001010010,
    17'b11111100101001000,
    17'b11111001111010111,
    17'b11110111000111101,
    17'b11110101000010100,
    17'b11110010001111011,
    17'b11101111010001111,
    17'b11101100000000000,
    17'b11101010110011010,
    17'b11101000101110001,
    17'b11100110100011111,
    17'b11100100111000011,
    17'b11100010101110001,
    17'b11100000100011111,
    17'b11011111001100110,
    17'b11011101001100110,
    17'b11011011010111000,
    17'b11011010101110001,
    17'b11011001101011100,
    17'b11011000101110001,
    17'b11011000101110001,
    17'b11011000010100100,
    17'b11010111100001010,
    17'b11010101110101110,
    17'b11010010101001000,
    17'b11010000000000000,
    17'b11001110011110110,
    17'b11001101000111101,
    17'b11001100000000000,
    17'b11000111001100110,
    17'b11000111001100110,
    17'b11000110111101100,
    17'b11000110101001000,
    17'b11000101010001111,
    17'b11000010100011111,
    17'b11000000111101100,
    17'b11000000100011111,
    17'b10111111110101110,
    17'b10111110111101100,
    17'b10111110001010010,
    17'b10111110010100100,
    17'b10111111111010111,
    17'b11000000111000011,
    17'b11000001110101110,
    17'b11000011010111000,
    17'b11000011001100110,
    17'b11000100001111011,
    17'b11000011110101110,
    17'b11000010101110001,
    17'b11000001100001010,
    17'b10111111110000101,
    17'b10111111011100001,
    17'b10111110010100100,
    17'b10111101110000101,
    17'b10111101100110011,
    17'b10111101010111000,
    17'b10111100110011010,
    17'b10111100111000011,
    17'b10111100101110001,
    17'b10111011010001111,
    17'b10111000111101100,
    17'b10110111100110011,
    17'b10110110101001000,
    17'b10110110011110110,
    17'b10110110011001101,
    17'b10110101000111101,
    17'b10110011010111000,
    17'b10110010110011010,
    17'b10110001010001111,
    17'b10101110010100100,
    17'b10101101010001111,
    17'b10101101100110011,
    17'b10101101110000101,
    17'b10101101110101110,
    17'b10101110011110110,
    17'b10101110001010010,
    17'b10101101100001010,
    17'b10101110000101001,
    17'b10101011110101110,
    17'b10101100001010010,
    17'b10101100000101001,
    17'b10101011100110011,
    17'b10101010000000000,
    17'b10101000111000011,
    17'b10101000111000011,
    17'b10101001010111000,
    17'b10101010111000011,
    17'b10101011000111101,
    17'b10101010100011111,
    17'b10101000111101100,
    17'b10101000011110110,
    17'b10100111000010100,
    17'b10100111010111000,
    17'b10100110010100100,
    17'b10100100111101100,
    17'b10100100100011111,
    17'b10100110001111011,
    17'b10100010101001000,
    17'b10100010001010010,
    17'b10100000000000000,
    17'b10011101111010111,
    17'b10011101010001111,
    17'b10011100011110110,
    17'b10011100111101100,
    17'b10011100111000011,
    17'b10011011101011100,
    17'b10011100001111011,
    17'b10011011110101110,
    17'b10011010110011010,
    17'b10011001101011100,
    17'b10011010110011010,
    17'b10011101001100110,
    17'b10011110111101100,
    17'b10011111110101110,
    17'b10100010101001000,
    17'b10100100010100100,
    17'b10100101000111101,
    17'b10100100110011010,
    17'b10100101000010100,
    17'b10100100011110110,
    17'b10100101001100110,
    17'b10100110011001101,
    17'b10101000011001101,
    17'b10101001110101110,
    17'b10101011010001111,
    17'b10101011100110011,
    17'b10101010101110001,
    17'b10100110101110001,
    17'b10100110111101100,
    17'b10100011000111101,
    17'b10100000100011111,
    17'b10011111101011100,
    17'b10011111011100001,
    17'b10011111100110011,
    17'b10011111000111101,
    17'b10011111010111000,
    17'b10100001000010100,
    17'b10100001000010100,
    17'b10100000101001000,
    17'b10011111111010111,
    17'b10100000101110001,
    17'b10100000101110001,
    17'b10011110101110001,
    17'b10011110111000011,
    17'b10011101101011100,
    17'b10011111000111101,
    17'b10011110000000000,
    17'b10011110001111011,
    17'b10011101011100001,
    17'b10011011110101110,
    17'b10011000001010010,
    17'b10010110010100100,
    17'b10010110110011010,
    17'b10011111000111101,
    17'b10011111110000101,
    17'b10011111001100110,
    17'b10011111100110011,
    17'b10100000111101100,
    17'b10100001110000101,
    17'b10100010101110001,
    17'b10100000111000011,
    17'b10011110111000011,
    17'b10011110010100100,
    17'b10011111010001111,
    17'b10011110111101100,
    17'b10011110011001101,
    17'b10011100000101001,
    17'b10011101000010100,
    17'b10011100011001101,
    17'b10011010110011010,
    17'b10011010001010010,
    17'b10011010100011111,
    17'b10011100000000000,
    17'b10011100010100100,
    17'b10011010101001000,
    17'b10011001011100001,
    17'b10011000110011010,
    17'b10010111110101110,
    17'b10011001001100110,
    17'b10011010001010010,
    17'b10011011110101110,
    17'b10011110011001101,
    17'b10100011100001010,
    17'b10100100000101001,
    17'b10101001100110011,
    17'b10110011001100110,
    17'b10110101100110011,
    17'b10111000111101100,
    17'b10111000110011010,
    17'b10111000000101001,
    17'b10110010110011010,
    17'b10101101110101110,
    17'b10101000010100100,
    17'b10100011100110011,
    17'b10011111010111000,
    17'b10011101111010111,
    17'b10011101100001010,
    17'b10011110001010010,
    17'b10011111011100001,
    17'b10100001010001111,
    17'b10100010110011010,
    17'b10100100100011111,
    17'b10100101100001010,
    17'b10100110000101001,
    17'b10100110100011111,
    17'b10101000000000000,
    17'b10101001100110011,
    17'b10101011101011100,
    17'b10110001111010111,
    17'b10110010101110001,
    17'b10110011100001010,
    17'b10110100000101001,
    17'b10110100011001101,
    17'b10110101010111000,
    17'b10110110010100100,
    17'b10110110111101100,
    17'b10110110100011111,
    17'b10110110000000000,
    17'b10110110001010010,
    17'b10110111010001111,
    17'b10111000101110001,
    17'b10111000011001101,
    17'b10110110101110001,
    17'b10110101000111101,
    17'b10110010100011111,
    17'b10110000011001101,
    17'b10101110100011111,
    17'b10101100111000011,
    17'b10101100100011111,
    17'b10101100111000011,
    17'b10101101100001010,
    17'b10101110111101100,
    17'b10110000101001000,
    17'b10110010001010010,
    17'b10110010101001000,
    17'b10110010101110001,
    17'b10110010101110001,
    17'b10110010011110110,
    17'b10110001100001010,
    17'b10110010000101001,
    17'b10110100001010010,
    17'b10110110001111011,
    17'b10111000100011111,
    17'b10111100000000000,
    17'b10111110011110110,
    17'b11000000111101100,
    17'b11000010101001000,
    17'b11000100101110001,
    17'b11000110001111011,
    17'b11000111000010100,
    17'b11000111100001010,
    17'b11000111100110011,
    17'b11000111001100110,
    17'b11000110011110110,
    17'b11000101111010111,
    17'b11000101010111000,
    17'b11000101011100001,
    17'b11000110000101001,
    17'b11000110101110001,
    17'b11001000000101001,
    17'b11001000111101100,
    17'b11001001100001010,
    17'b11001010011001101,
    17'b11001010110011010,
    17'b11001010111101100,
    17'b11001010001111011,
    17'b11001001101011100,
    17'b11001010010100100,
    17'b11001010101110001,
    17'b11001010111000011,
    17'b11001011111010111,
    17'b11001101011100001,
    17'b11001110101110001,
    17'b11010111100001010,
    17'b11011011110101110,
    17'b11011111111010111,
    17'b11100010111101100,
    17'b11100100000101001,
    17'b11100101010001111,
    17'b11100110001010010,
    17'b11100110001010010,
    17'b11100101001100110,
    17'b11100011101011100,
    17'b11100011100110011,
    17'b11100010111000011,
    17'b11100011000010100,
    17'b11100011010001111,
    17'b11100011011100001,
    17'b11100011011100001,
    17'b11100011100001010,
    17'b11100011100110011,
    17'b11100011101011100,
    17'b11100100000000000,
    17'b11100100001010010,
    17'b11100011100110011,
    17'b11100010111000011,
    17'b11100001111010111,
    17'b11100001110101110,
    17'b11100010001010010,
    17'b11100011010111000,
    17'b11100100000000000,
    17'b11100101000010100,
    17'b11100101110101110,
    17'b11100110011110110,
    17'b11100111000010100,
    17'b11100111110101110,
    17'b11101000011001101,
    17'b11101001010111000,
    17'b11101001010111000,
    17'b11101001010111000,
    17'b11101001100001010,
    17'b11101010011001101,
    17'b11101011110101110,
    17'b11101101000111101,
    17'b11101110001010010,
    17'b11101011000111101,
    17'b11101010011001101,
    17'b11101010010100100,
    17'b11101010001111011,
    17'b11101001010111000,
    17'b11100111111010111,
    17'b11100111001100110,
    17'b11100110101001000,
    17'b11100101111010111,
    17'b11100101110000101,
    17'b11100110001010010,
    17'b11101000001111011,
    17'b11101000000000000,
    17'b11101000101110001,
    17'b11101001100110011,
    17'b11101001010001111,
    17'b11101000111000011,
    17'b11101010000000000,
    17'b11101100101001000,
    17'b11101110101001000,
    17'b11110000001010010,
    17'b11110010010100100,
    17'b11110010011001101,
    17'b11110011000010100,
    17'b11110100011110110,
    17'b11110110101110001,
    17'b11110110111000011,
    17'b11110110111101100,
    17'b11110111001100110,
    17'b11110011011100001,
    17'b11101111110000101,
    17'b11101111110101110,
    17'b11110100000000000,
    17'b11110110110011010,
    17'b11111001101011100,
    17'b11111011100110011,
    17'b11111011100001010,
    17'b11111000001111011,
    17'b11110110111000011,
    17'b11110000011110110,
    17'b11110010001010010,
    17'b11110011110101110,
    17'b11110110011110110,
    17'b11110111000111101,
    17'b11111000111000011,
    17'b11111010011001101,
    17'b11111011010111000,
    17'b11111101010111000,
    17'b11111110100011111,
    17'b11111110101001000,
    17'b11111111010111000,
    17'b11111111011100001,
    17'b11111111100110011,
    17'b11111111101011100,
    17'b11111111100001010,
    17'b11111111000111101,
    17'b11111110110011010,
    17'b11111111001100110,
    17'b11111110000000000,
    17'b11111110000101001,
    17'b11111101100110011,
    17'b11111110011110110,
    17'b11111111111010111,
    17'b00000001100001010,
    17'b00000001000010100,
    17'b00000001111010111,
    17'b00000010110011010,
    17'b00000010101110001,
    17'b00000100010100100,
    17'b00000101010111000,
    17'b00000100001111011,
    17'b00000111001100110,
    17'b00010111101011100,
    17'b00001100101001000,
    17'b00001100101110001,
    17'b00001100001010010,
    17'b00001100101110001,
    17'b00001011010111000,
    17'b00001001010111000,
    17'b00001000001010010,
    17'b00001000110011010,
    17'b00001010001010010,
    17'b00001101001100110,
    17'b00001110000000000,
    17'b00010001100110011,
    17'b00010010001111011,
    17'b00010010000000000,
    17'b00010001100110011,
    17'b00010000000101001,
    17'b00001111000010100,
    17'b00001110001010010,
    17'b00001110100011111,
    17'b00001110001111011,
    17'b00001110011001101,
    17'b00001110110011010,
    17'b00001111011100001,
    17'b00010000001111011,
    17'b00010010011110110,
    17'b00010010010100100,
    17'b00001110010100100,
    17'b00001101100110011,
    17'b00010001000111101,
    17'b00010100110011010,
    17'b00010010101110001,
    17'b00010000011001101,
    17'b00001111110101110,
    17'b00010001111010111,
    17'b00001111001100110,
    17'b00001111100110011,
    17'b00010001011100001,
    17'b00010111100001010,
    17'b00001110000000000,
    17'b00001100111000011,
    17'b00001110000101001,
    17'b00010011101011100,
    17'b00010011110101110,
    17'b00001100000101001,
    17'b00001111011100001,
    17'b00010101110101110,
    17'b00001101010001111,
    17'b00010100011001101,
    17'b00001101010111000,
    17'b00001101010001111,
    17'b00010011100001010,
    17'b00001110101001000,
    17'b00001011110000101,
    17'b00010111010111000,
    17'b00011101000010100,
    17'b00001110001111011,
    17'b00100000001111011,
    17'b00011110101110001,
    17'b00011100110011010,
    17'b00100001000111101,
    17'b00100000000101001,
    17'b00100010101110001,
    17'b00001011001100110,
    17'b00001011000010100,
    17'b00001010000000000,
    17'b00000111010001111,
    17'b11110111010111000,
    17'b11111111100110011,
    17'b00000010100011111,
    17'b00001000001010010,
    17'b00001011000111101,
    17'b00001010100011111,
    17'b00000111110101110,
    17'b00000110011001101,
    17'b00000101001100110,
    17'b00000100100011111,
    17'b00000100011001101,
    17'b00000100000101001,
    17'b00000011011100001,
    17'b00000010111101100,
    17'b00000010001111011,
    17'b00000001010001111,
    17'b11111110101001000,
    17'b11111011100001010,
    17'b11111010000101001,
    17'b11111001001100110,
    17'b11111000001010010,
    17'b11111001011100001,
    17'b11110111101011100,
    17'b11110111000111101,
    17'b11110110001010010,
    17'b11110101001100110,
    17'b11110100011110110,
    17'b11110010111000011,
    17'b11110001100001010,
    17'b11110000000000000,
    17'b11101110111101100,
    17'b11101110000101001,
    17'b11101100111000011,
    17'b11101100001111011,
    17'b11101011100110011,
    17'b11101010110011010,
    17'b11100111000111101,
    17'b11100110011110110,
    17'b11100101101011100,
    17'b11100100110011010,
    17'b11100100011001101,
    17'b11100100000000000,
    17'b11100011111010111,
    17'b11100010101001000,
    17'b11100001000111101,
    17'b11011101000111101,
    17'b11011010010100100,
    17'b11011001000111101,
    17'b11011000001111011,
    17'b11010111011100001,
    17'b11010110011001101,
    17'b11010101001100110,
    17'b11010011110000101,
    17'b11010010011110110,
    17'b11010001111010111,
    17'b11010001000111101,
    17'b11010000010100100,
    17'b11010000000101001,
    17'b11010000101001000,
    17'b11010001010111000,
    17'b11010101010111000,
    17'b11010100010100100,
    17'b11001110011110110,
    17'b11010000010100100,
    17'b11001110110011010,
    17'b11000111101011100,
    17'b11000100000000000,
    17'b10111010111101100,
    17'b10111010100011111,
    17'b10111011000010100,
    17'b10111011100001010,
    17'b10111011011100001,
    17'b10111010101001000,
    17'b10111001110000101,
    17'b10111001110000101,
    17'b10111011111010111,
    17'b10111010010100100,
    17'b10111000000000000,
    17'b10111000011110110,
    17'b10110101110101110,
    17'b10110100101110001,
    17'b10110100110011010,
    17'b10110100011001101,
    17'b10110100101110001,
    17'b10110110100011111,
    17'b10110111110101110,
    17'b10110110001111011,
    17'b10110101110101110,
    17'b10110111010111000,
    17'b10110101100110011,
    17'b10110000101001000,
    17'b10110001101011100,
    17'b10101110001010010,
    17'b10100110111101100,
    17'b10100101000010100,
    17'b10100100101110001,
    17'b10100001100001010,
    17'b10100011001100110,
    17'b10100011111010111,
    17'b10100001110000101,
    17'b10100000010100100,
    17'b10011111010001111,
    17'b10011101011100001,
    17'b10011011110000101,
    17'b10011100011001101,
    17'b10011100111101100,
    17'b10011100111101100,
    17'b10011100111101100,
    17'b10011100011001101,
    17'b10011100101001000,
    17'b10011101110101110,
    17'b10011101111010111,
    17'b10011110001010010,
    17'b10011101010111000,
    17'b10011100111000011,
    17'b10011011110101110,
    17'b10011011000111101,
    17'b10011010000101001,
    17'b10011010100011111,
    17'b10011010000101001,
    17'b10011011110000101,
    17'b10011101011100001,
    17'b10100000101110001,
    17'b10100000101110001,
    17'b10011111110000101,
    17'b10011111011100001,
    17'b10011110101001000,
    17'b10011110000000000,
    17'b10011100111000011,
    17'b10011011101011100,
    17'b10011010011110110,
    17'b10011001101011100,
    17'b10011001111010111,
    17'b10011010011110110,
    17'b10011011111010111,
    17'b10011100010100100,
    17'b10011101101011100,
    17'b10011110111000011,
    17'b10011111101011100,
    17'b10100000010100100,
    17'b10011111000010100,
    17'b10011110111000011,
    17'b10011111000111101,
    17'b10011111010111000,
    17'b10011101111010111,
    17'b10011101100001010,
    17'b10011011111010111,
    17'b10011101001100110,
    17'b10011110001010010,
    17'b10011110111101100,
    17'b10011111010111000,
    17'b10011111101011100,
    17'b10100001000010100,
    17'b10100010001111011,
    17'b10100011001100110,
    17'b10100100001111011,
    17'b10100100000101001,
    17'b10100100101001000,
    17'b10100100011110110,
    17'b10100100111000011,
    17'b10100101110000101,
    17'b10100111010001111,
    17'b10101000001111011,
    17'b10101000011110110,
    17'b10110010011110110,
    17'b10111111010001111,
    17'b10111000110011010,
    17'b10110101101011100,
    17'b10110010001111011,
    17'b10110000001010010,
    17'b10101110111101100,
    17'b10101001100001010,
    17'b10100100000101001,
    17'b10100010000000000,
    17'b10011111000111101,
    17'b10011110110011010,
    17'b10011111100110011,
    17'b10100001100110011,
    17'b10100100011001101,
    17'b10101100000101001,
    17'b10101101010111000,
    17'b10100110111000011,
    17'b10100011010111000,
    17'b10011010111101100,
    17'b10011100000000000,
    17'b10011110111101100,
    17'b10100010111101100,
    17'b10100110000101001,
    17'b10101001101011100,
    17'b10101010110011010,
    17'b10101010111000011,
    17'b10101001000111101,
    17'b10100111000111101,
    17'b10100101000010100,
    17'b10100011000010100,
    17'b10100000010100100,
    17'b10011100111000011,
    17'b10011010101001000,
    17'b10011001011100001,
    17'b10011011000010100,
    17'b10011101000010100,
    17'b10011101000010100,
    17'b10011100001111011,
    17'b10011011010001111,
    17'b10011101000010100,
    17'b10011110100011111,
    17'b10011101000111101,
    17'b10011100001010010,
    17'b10011101110000101,
    17'b10011010101110001,
    17'b10100011000010100,
    17'b10101000011110110,
    17'b10101000100011111,
    17'b10101000000101001,
    17'b10101000111101100,
    17'b10101001111010111,
    17'b10101011011100001,
    17'b10101100001111011,
    17'b10101101101011100,
    17'b10101110001010010,
    17'b10101101100110011,
    17'b10101100000000000,
    17'b10101010011110110,
    17'b10101000000101001,
    17'b10100101100001010,
    17'b10100001110101110,
    17'b10011111011100001,
    17'b10011101100001010,
    17'b10011011011100001,
    17'b10011010011110110,
    17'b10011010010100100,
    17'b10011010111000011,
    17'b10011100111000011,
    17'b10100110000000000,
    17'b10100111110101110,
    17'b10101010001111011,
    17'b10101011110000101,
    17'b10101100111000011,
    17'b10101110000101001,
    17'b10101110110011010,
    17'b10101111000111101,
    17'b10101111010001111,
    17'b10110000000000000,
    17'b10101111000111101,
    17'b10101110111101100,
    17'b10101110001010010,
    17'b10101110000101001,
    17'b10101101101011100,
    17'b10101100100011111,
    17'b10101010010100100,
    17'b10101000011110110,
    17'b10100101110101110,
    17'b10100100001010010,
    17'b10100010011001101,
    17'b10100010000101001,
    17'b10100010001111011,
    17'b10100010011001101,
    17'b10100010100011111,
    17'b10100011110101110,
    17'b10100101011100001,
    17'b10101100101110001,
    17'b10101100101001000,
    17'b10101011100001010,
    17'b10101000010100100,
    17'b10101000111101100,
    17'b10101010010100100,
    17'b10101011110000101,
    17'b10011000011001101,
    17'b10011000111000011,
    17'b10100001110101110,
    17'b10100110001010010,
    17'b10100111100001010,
    17'b10101110001010010,
    17'b10110001110101110,
    17'b10110010011110110,
    17'b10110011111010111,
    17'b10110100101110001,
    17'b10110111010001111,
    17'b10110110011001101,
    17'b10110100001111011,
    17'b10110101100110011,
    17'b10110100110011010,
    17'b10110001011100001,
    17'b10110000010100100,
    17'b10101111100001010,
    17'b10101110010100100,
    17'b10101101001100110,
    17'b10101100010100100,
    17'b10101011000111101,
    17'b10101001101011100,
    17'b10101001010001111,
    17'b10101010001111011,
    17'b10101100001010010,
    17'b10101101111010111,
    17'b10110010011001101,
    17'b10110011000010100,
    17'b10110011001100110,
    17'b10110100011110110,
    17'b10110110011110110,
    17'b10111000011001101,
    17'b10111010010100100,
    17'b10111100001111011,
    17'b10111110111000011,
    17'b11000001101011100,
    17'b11000011100110011,
    17'b11000100010100100,
    17'b11000101000010100,
    17'b11000101001100110,
    17'b11000100111101100,
    17'b11000100011001101,
    17'b11000011100110011,
    17'b11000011010111000,
    17'b11000010101110001,
    17'b11000000110011010,
    17'b10111101010001111,
    17'b10111011101011100,
    17'b10111011000111101,
    17'b10111010101001000,
    17'b10111010000101001,
    17'b10111001010111000,
    17'b10111000111101100,
    17'b10111001111010111,
    17'b10111011011100001,
    17'b10111100000101001,
    17'b10111011001100110,
    17'b10111010100011111,
    17'b10111011001100110,
    17'b10111011010001111,
    17'b10111011010001111,
    17'b10111100011001101,
    17'b10111101111010111,
    17'b10111111010001111,
    17'b11000001101011100,
    17'b11000010000101001,
    17'b11000011111010111,
    17'b11000010100011111,
    17'b11000110101110001,
    17'b11001111010111000,
    17'b11010010011110110,
    17'b11010110001111011,
    17'b11011010011001101,
    17'b11011001100001010,
    17'b11010111010001111,
    17'b11010101110101110,
    17'b11010100100011111,
    17'b11010100110011010,
    17'b11010100111101100,
    17'b11010101010001111,
    17'b11010101111010111,
    17'b11010110000000000,
    17'b11010110011110110,
    17'b11010111010111000,
    17'b11011000010100100,
    17'b11011001000010100,
    17'b11011010000101001,
    17'b11011011100110011,
    17'b11011100111101100,
    17'b11011101101011100,
    17'b11011110000000000,
    17'b11011110010100100,
    17'b11011110111101100,
    17'b11100000001010010,
    17'b11100001110101110,
    17'b11100100000000000,
    17'b11100101110101110,
    17'b11100111100110011,
    17'b11101001000010100,
    17'b11101011100110011,
    17'b11101101101011100,
    17'b11101111100110011,
    17'b11110000111101100,
    17'b11110010101110001,
    17'b11110011111010111,
    17'b11110100111101100,
    17'b11111010010100100,
    17'b11111011111010111,
    17'b11111100011110110,
    17'b11111101110000101,
    17'b11111111011100001,
    17'b00000000001010010,
    17'b00000001000111101,
    17'b00000010011001101,
    17'b00000100011001101,
    17'b00000110010100100,
    17'b00000110111000011,
    17'b00001001111010111,
    17'b00001001111010111,
    17'b00001010011001101,
    17'b00001100000101001,
    17'b00001110111101100,
    17'b00001111100110011,
    17'b00010010000000000,
    17'b00010001110101110,
    17'b00010010001111011,
    17'b00010010111101100,
    17'b00010100011001101,
    17'b00010110001111011,
    17'b00010111110101110,
    17'b00011001100001010,
    17'b00011011001100110,
    17'b00011100011110110,
    17'b00011101010111000,
    17'b00011110101001000,
    17'b00011111110101110,
    17'b00100000101001000,
    17'b00100001101011100,
    17'b00100011010001111,
    17'b00100100100011111,
    17'b00100101101011100,
    17'b00100101110101110,
    17'b00100110000000000,
    17'b00100101001100110,
    17'b00100101000010100,
    17'b00100101011100001,
    17'b00100101110000101,
    17'b00100110001010010,
    17'b00100110010100100,
    17'b00100110110011010,
    17'b00100111100001010,
    17'b00101001001100110,
    17'b00101100001111011,
    17'b00101110111000011,
    17'b00110001010111000,
    17'b00110010111000011,
    17'b00110010101001000,
    17'b00110010101110001,
    17'b00110011000111101,
    17'b00110010101110001,
    17'b00110010101110001,
    17'b00110010111101100,
    17'b00110010000101001,
    17'b00101111111010111,
    17'b00101110100011111,
    17'b00101101101011100,
    17'b00101011101011100,
    17'b00101011000111101,
    17'b00101011010111000,
    17'b00101011001100110,
    17'b00101010010100100,
    17'b00101001000010100
};

parameter logic signed [`GYRO_WIDTH-1:0] WX_TEST_VECTOR[`NUM_ELEMENTS] = {
    22'b1111110001111010111000,
    22'b1111110001110000101001,
    22'b1111110001011100001010,
    22'b1111110001000111101100,
    22'b1111110000011110101110,
    22'b1111101111010111000011,
    22'b1111101110011001100110,
    22'b1111101101000111101100,
    22'b1111101011101011100001,
    22'b1111101001011100001010,
    22'b1111100111100001010010,
    22'b1111100101011100001010,
    22'b1111100011010111000011,
    22'b1111100000101000111101,
    22'b1111011110111000010100,
    22'b1111011101100110011010,
    22'b1111011100111101011100,
    22'b1111011100110011001101,
    22'b1111011101000111101100,
    22'b1111011101111010111000,
    22'b1111011111000010100100,
    22'b1111100000111101011100,
    22'b1111100010011001100110,
    22'b1111100011101011100001,
    22'b1111100100110011001101,
    22'b1111100101111010111000,
    22'b1111100110011001100110,
    22'b1111100110101110000101,
    22'b1111100110101110000101,
    22'b1111100110001111010111,
    22'b1111100101100110011010,
    22'b1111100100110011001101,
    22'b1111100011010111000011,
    22'b1111100010011001100110,
    22'b1111100001000111101100,
    22'b1111100000010100011111,
    22'b1111100000101000111101,
    22'b1111100001011100001010,
    22'b1111100010101110000101,
    22'b1111100100000000000000,
    22'b1111100100110011001101,
    22'b1111100100110011001101,
    22'b1111100100011110101110,
    22'b1111100100011110101110,
    22'b1111100100111101011100,
    22'b1111100101111010111000,
    22'b1111100111010111000011,
    22'b1111101000110011001101,
    22'b1111101011000010100100,
    22'b1111101100110011001101,
    22'b1111101110101110000101,
    22'b1111110000101000111101,
    22'b1111110011010111000011,
    22'b1111110101011100001010,
    22'b1111110111101011100001,
    22'b1111111010100011110110,
    22'b1111111100101000111101,
    22'b1111111110001111010111,
    22'b1111111111001100110011,
    22'b0000000000000000000000,
    22'b0000000000000000000000,
    22'b1111111111110101110001,
    22'b1111111111100001010010,
    22'b1111111110011001100110,
    22'b1111111100111101011100,
    22'b1111111011110101110001,
    22'b1111111011100001010010,
    22'b1111111100101000111101,
    22'b1111111110101110000101,
    22'b0000000001111010111000,
    22'b0000000101111010111000,
    22'b0000001011001100110011,
    22'b0000001101111010111000,
    22'b0000001111000010100100,
    22'b0000001110100011110110,
    22'b0000001001111010111000,
    22'b0000000011001100110011,
    22'b1111111011101011100001,
    22'b1111111100111101011100,
    22'b0000000001010001111011,
    22'b0000001011110101110001,
    22'b0000011100101000111101,
    22'b0000110101010001111011,
    22'b0001000100011110101110,
    22'b0001001010101110000101,
    22'b0000111110011001100110,
    22'b0000101000111101011100,
    22'b0000010000001010001111,
    22'b1111111011000010100100,
    22'b1111101001011100001010,
    22'b1111100101110000101001,
    22'b1111101000001010001111,
    22'b1111101110000101001000,
    22'b1111110111101011100001,
    22'b1111111110000101001000,
    22'b0000000011001100110011,
    22'b0000000111010111000011,
    22'b0000001011101011100001,
    22'b0000001110000101001000,
    22'b0000001111110101110001,
    22'b0000010010001111010111,
    22'b0000010100010100011111,
    22'b0000010110000101001000,
    22'b0000010110111000010100,
    22'b0000010110101110000101,
    22'b0000010110001111010111,
    22'b0000010100101000111101,
    22'b0000010001111010111000,
    22'b0000001110101110000101,
    22'b0000001010101110000101,
    22'b0000000110100011110110,
    22'b0000000001010001111011,
    22'b1111111110100011110110,
    22'b1111111101010001111011,
    22'b1111111101011100001010,
    22'b1111111111000010100100,
    22'b0000000000101000111101,
    22'b0000000010100011110110,
    22'b0000000100010100011111,
    22'b0000000101011100001010,
    22'b0000000101010001111011,
    22'b0000000011100001010010,
    22'b1111111100101000111101,
    22'b1111111000111101011100,
    22'b1111111000001010001111,
    22'b1111110111001100110011,
    22'b1111110101111010111000,
    22'b1111110101000111101100,
    22'b1111110100101000111101,
    22'b1111110011110101110001,
    22'b1111110011100001010010,
    22'b1111110011110101110001,
    22'b1111110101010001111011,
    22'b1111110111000010100100,
    22'b1111111000010100011111,
    22'b1111111001110000101001,
    22'b1111111100001010001111,
    22'b1111111101011100001010,
    22'b1111111101100110011010,
    22'b1111111110111000010100,
    22'b1111111111010111000011,
    22'b1111111101110000101001,
    22'b1111111100010100011111,
    22'b1111111100001010001111,
    22'b1111111100000000000000,
    22'b1111111100110011001101,
    22'b1111111101011100001010,
    22'b1111111001011100001010,
    22'b1111110100111101011100,
    22'b1111110001111010111000,
    22'b1111101111101011100001,
    22'b1111101101111010111000,
    22'b1111101011110101110001,
    22'b1111101001111010111000,
    22'b1111101000011110101110,
    22'b1111101001000111101100,
    22'b1111101000000000000000,
    22'b1111100111001100110011,
    22'b1111100110001111010111,
    22'b1111100101011100001010,
    22'b1111100011110101110001,
    22'b1111100010101110000101,
    22'b1111100001011100001010,
    22'b1111100000110011001101,
    22'b1111100000011110101110,
    22'b1111100001100110011010,
    22'b1111100100000000000000,
    22'b1111100111001100110011,
    22'b1111101010011001100110,
    22'b1111101100101000111101,
    22'b1111101110101110000101,
    22'b1111110000010100011111,
    22'b1111110001011100001010,
    22'b1111110001011100001010,
    22'b1111110000101000111101,
    22'b1111101111101011100001,
    22'b1111101110011001100110,
    22'b1111101100101000111101,
    22'b1111101010101110000101,
    22'b1111101010101110000101,
    22'b1111101011001100110011,
    22'b1111101011100001010010,
    22'b1111101000110011001101,
    22'b1111100111010111000011,
    22'b1111100101010001111011,
    22'b1111100100010100011111,
    22'b1111100110000101001000,
    22'b1111101011100001010010,
    22'b1111110110101110000101,
    22'b1111111010100011110110,
    22'b1111111110101110000101,
    22'b0000000010001111010111,
    22'b0000000010011001100110,
    22'b1111111111101011100001,
    22'b1111111100110011001101,
    22'b1111111010011001100110,
    22'b1111111000011110101110,
    22'b1111110111100001010010,
    22'b1111110110100011110110,
    22'b1111110100000000000000,
    22'b1111101110101110000101,
    22'b1111101110111000010100,
    22'b1111101111000010100100,
    22'b1111101000011110101110,
    22'b1111100001000111101100,
    22'b1111100001011100001010,
    22'b1111011111000010100100,
    22'b1111011101000111101100,
    22'b1111100010000101001000,
    22'b1111100110000101001000,
    22'b1111101001011100001010,
    22'b1111101101100110011010,
    22'b1111110010001111010111,
    22'b1111111000110011001101,
    22'b1111111111001100110011,
    22'b0000000110111000010100,
    22'b0000001110111000010100,
    22'b0000010111000010100100,
    22'b0000011010101110000101,
    22'b0000011011110101110001,
    22'b0000011010000101001000,
    22'b0000010010101110000101,
    22'b0000001010111000010100,
    22'b0000000001111010111000,
    22'b1111111001000111101100,
    22'b1111110000110011001101,
    22'b1111100111110101110001,
    22'b1111100010111000010100,
    22'b1111011111110101110001,
    22'b1111011110000101001000,
    22'b1111011101011100001010,
    22'b1111011101111010111000,
    22'b1111011110100011110110,
    22'b1111011111010111000011,
    22'b1111100000111101011100,
    22'b1111100010100011110110,
    22'b1111100100110011001101,
    22'b1111101000010100011111,
    22'b1111101011010111000011,
    22'b1111101110101110000101,
    22'b1111110010011001100110,
    22'b1111110111101011100001,
    22'b1111111011100001010010,
    22'b1111111111100001010010,
    22'b0000000010011001100110,
    22'b1111111000010100011111,
    22'b1111101011110101110001,
    22'b1111101001110000101001,
    22'b1111101010000101001000,
    22'b1111100100001010001111,
    22'b1111011111000010100100,
    22'b1111100001100110011010,
    22'b1111011100000000000000,
    22'b1111011010101110000101,
    22'b1111011111101011100001,
    22'b1111101001010001111011,
    22'b1111110100110011001101,
    22'b1111111011000010100100,
    22'b0000000000000000000000,
    22'b0000000010000101001000,
    22'b0000000011010111000011,
    22'b0000000010011001100110,
    22'b0000000000111101011100,
    22'b0000000001100110011010,
    22'b0000000001011100001010,
    22'b0000000001000111101100,
    22'b0000000000110011001101,
    22'b0000000000110011001101,
    22'b0000000000101000111101,
    22'b0000000001000111101100,
    22'b0000000000110011001101,
    22'b1111111111110101110001,
    22'b0000000000010100011111,
    22'b0000000000101000111101,
    22'b0000000000111101011100,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000000101000111101,
    22'b0000000000111101011100,
    22'b0000000001000111101100,
    22'b0000000000101000111101,
    22'b1111111111001100110011,
    22'b1111111101111010111000,
    22'b1111111111010111000011,
    22'b0000000001011100001010,
    22'b0000000010101110000101,
    22'b0000000011101011100001,
    22'b0000000010001111010111,
    22'b0000000001100110011010,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001110000101001,
    22'b0000000001100110011010,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001010001111011,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001000111101100,
    22'b0000000000111101011100,
    22'b0000000000110011001101,
    22'b0000000000101000111101,
    22'b0000000000010100011111,
    22'b1111111111110101110001,
    22'b1111111111001100110011,
    22'b1111111111110101110001,
    22'b0000000001010001111011,
    22'b0000000011001100110011,
    22'b0000000010011001100110,
    22'b0000000001111010111000,
    22'b0000000001111010111000,
    22'b0000000001110000101001,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001000111101100,
    22'b0000000001011100001010,
    22'b0000000001100110011010,
    22'b0000000001100110011010,
    22'b0000000001100110011010,
    22'b0000000001010001111011,
    22'b0000000000110011001101,
    22'b0000000000110011001101,
    22'b0000000001000111101100,
    22'b0000000001010001111011,
    22'b0000000001100110011010,
    22'b0000000001111010111000,
    22'b0000000001110000101001,
    22'b0000000001100110011010,
    22'b0000000001011100001010,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000000111101011100,
    22'b1111111010111000010100,
    22'b1111101111001100110011,
    22'b1111100000001010001111,
    22'b1111100000110011001101,
    22'b1111100010111000010100,
    22'b1111101000010100011111,
    22'b1111101101111010111000,
    22'b1111110110101110000101,
    22'b1111111110000101001000,
    22'b0000000100110011001101,
    22'b0000000111001100110011,
    22'b0000000110111000010100,
    22'b0000000000010100011111,
    22'b1111111110000101001000,
    22'b1111111000110011001101,
    22'b1111101100001010001111,
    22'b1111000011010111000011,
    22'b1110011000001010001111,
    22'b1110100111001100110011,
    22'b1110110101100110011010,
    22'b1111010101111010111000,
    22'b1111111100000000000000,
    22'b0000101100010100011111,
    22'b0001010001011100001010,
    22'b0001100100110011001101,
    22'b0001101110001111010111,
    22'b0001001011101011100001,
    22'b0000101011101011100001,
    22'b0000011110001111010111,
    22'b0000011110101110000101,
    22'b0000010111001100110011,
    22'b0000010011101011100001,
    22'b0000001101010001111011,
    22'b0000001001000111101100,
    22'b0000000101010001111011,
    22'b0000000010011001100110,
    22'b1111111110011001100110,
    22'b1111111010001111010111,
    22'b1111110001111010111000,
    22'b1111101101100110011010,
    22'b1111101000001010001111,
    22'b1111100000000000000000,
    22'b1111011011001100110011,
    22'b1111011001110000101001,
    22'b1111011110000101001000,
    22'b1111101101000111101100,
    22'b1111111101111010111000,
    22'b0000010000011110101110,
    22'b0000100001111010111000,
    22'b0000101111101011100001,
    22'b0000111000000000000000,
    22'b0000011110000101001000,
    22'b0000010100000000000000,
    22'b0000010011100001010010,
    22'b0000001100010100011111,
    22'b0000000010100011110110,
    22'b0000000010101110000101,
    22'b0000000011001100110011,
    22'b0000000010101110000101,
    22'b0000000011000010100100,
    22'b0000000010011001100110,
    22'b0000000010100011110110,
    22'b1111111111001100110011,
    22'b1111111001010001111011,
    22'b1111110100101000111101,
    22'b1111110000111101011100,
    22'b1111101110100011110110,
    22'b1111101111101011100001,
    22'b1111110010111000010100,
    22'b1111110111110101110001,
    22'b0000000000010100011111,
    22'b0000000111001100110011,
    22'b0000001101100110011010,
    22'b0000010011001100110011,
    22'b0000010111101011100001,
    22'b0000001101110000101001,
    22'b0000001011101011100001,
    22'b0000001000101000111101,
    22'b0000000101100110011010,
    22'b0000000100001010001111,
    22'b0000000011001100110011,
    22'b0000000010100011110110,
    22'b0000000010001111010111,
    22'b0000000001110000101001,
    22'b0000000001100110011010,
    22'b0000000001011100001010,
    22'b0000000000110011001101,
    22'b1111111110100011110110,
    22'b1111111101100110011010,
    22'b1111111100111101011100,
    22'b1111111100011110101110,
    22'b1111111100101000111101,
    22'b1111111101011100001010,
    22'b1111111110101110000101,
    22'b0000000001010001111011,
    22'b0000000011110101110001,
    22'b0000000110011001100110,
    22'b0000001000010100011111,
    22'b0000000101011100001010,
    22'b0000000100010100011111,
    22'b0000000011010111000011,
    22'b0000000010101110000101,
    22'b0000000010001111010111,
    22'b0000000001110000101001,
    22'b0000000001100110011010,
    22'b0000000001111010111000,
    22'b0000000010001111010111,
    22'b0000000010011001100110,
    22'b0000000010111000010100,
    22'b0000000010100011110110,
    22'b0000000100010100011111,
    22'b0000000100101000111101,
    22'b1111111100000000000000,
    22'b1111110001011100001010,
    22'b1111101101011100001010,
    22'b1111110100011110101110,
    22'b1111110101010001111011,
    22'b1111111011010111000011,
    22'b0000001011101011100001,
    22'b0000011011110101110001,
    22'b0000100011110101110001,
    22'b0000011111010111000011,
    22'b0000101110101110000101,
    22'b0001000110100011110110,
    22'b0001001010101110000101,
    22'b0001000111110101110001,
    22'b0001001000011110101110,
    22'b0001010100010100011111,
    22'b0001011000101000111101,
    22'b0001001011100001010010,
    22'b0000111100101000111101,
    22'b0000110010000101001000,
    22'b0000110011001100110011,
    22'b0000111001011100001010,
    22'b0001000011010111000011,
    22'b0001010010011001100110,
    22'b0001010111110101110001,
    22'b0001010111010111000011,
    22'b0001010100101000111101,
    22'b0001001101110000101001,
    22'b0001000111100001010010,
    22'b0001000001111010111000,
    22'b0000111101110000101001,
    22'b0000111010111000010100,
    22'b0000110111010111000011,
    22'b0000110100011110101110,
    22'b0000110001010001111011,
    22'b0000101100101000111101,
    22'b0000100111000010100100,
    22'b0000100101010001111011,
    22'b0000100100010100011111,
    22'b0000100010111000010100,
    22'b0000100001010001111011,
    22'b0000011111101011100001,
    22'b0000011101011100001010,
    22'b0000011011010111000011,
    22'b0000011010000101001000,
    22'b0000011001111010111000,
    22'b0000011000110011001101,
    22'b0000010111000010100100,
    22'b0000010011000010100100,
    22'b0000010011100001010010,
    22'b0000010110011001100110,
    22'b0000010111100001010010,
    22'b0000010110111000010100,
    22'b0000010100111101011100,
    22'b0000010100101000111101,
    22'b0000010010101110000101,
    22'b0000001101110000101001,
    22'b0000001001110000101001,
    22'b0000000101100110011010,
    22'b0000000010100011110110,
    22'b0000000010100011110110,
    22'b0000000101010001111011,
    22'b0000001000110011001101,
    22'b0000001101000111101100,
    22'b0000001111110101110001,
    22'b0000010001111010111000,
    22'b0000010100001010001111,
    22'b0000010101111010111000,
    22'b0000011000101000111101,
    22'b0000011010000101001000,
    22'b0000011001000111101100,
    22'b0000011001011100001010,
    22'b0000011001100110011010,
    22'b0000001010111000010100,
    22'b1111111001000111101100,
    22'b1111111011001100110011,
    22'b0000000001000111101100,
    22'b0000000101010001111011,
    22'b0000001100011110101110,
    22'b0000010011101011100001,
    22'b0000011000111101011100,
    22'b0000100010100011110110,
    22'b0000110001000111101100,
    22'b0000111010111000010100,
    22'b0000111000010100011111,
    22'b0000111000001010001111,
    22'b0000110100110011001101,
    22'b0000100101011100001010,
    22'b0000101100011110101110,
    22'b0000101010011001100110,
    22'b0000110000010100011111,
    22'b0001000001000111101100,
    22'b0001000111001100110011,
    22'b0001000101111010111000,
    22'b0000111111010111000011,
    22'b0000111110000101001000,
    22'b0000111101100110011010,
    22'b0000111101111010111000,
    22'b0000111001111010111000,
    22'b0000111000110011001101,
    22'b0000110011110101110001,
    22'b0000101101011100001010,
    22'b0000100010001111010111,
    22'b0000011000110011001101,
    22'b0000000110001111010111,
    22'b1111101110000101001000,
    22'b1111001000010100011111,
    22'b1110110010111000010100,
    22'b1110100011101011100001,
    22'b1110011110001111010111,
    22'b1110100011110101110001,
    22'b1111001010101110000101,
    22'b0000100000010100011111,
    22'b0001000101011100001010,
    22'b0000110100010100011111,
    22'b0000011011010111000011,
    22'b0000001011110101110001,
    22'b0000010011000010100100,
    22'b0000111110101110000101,
    22'b0001011101111010111000,
    22'b0001100100010100011111,
    22'b0001010101100110011010,
    22'b0000111111000010100100,
    22'b0000100110100011110110,
    22'b0000100011101011100001,
    22'b0000100010111000010100,
    22'b0000100111100001010010,
    22'b0000111010100011110110,
    22'b0001000110100011110110,
    22'b0001001010000101001000,
    22'b0001001010111000010100,
    22'b0001001111010111000011,
    22'b0001011000010100011111,
    22'b0001011110001111010111,
    22'b0001100100001010001111,
    22'b0001101000111101011100,
    22'b0001101110011001100110,
    22'b0001110010001111010111,
    22'b0001110110100011110110,
    22'b0001111001111010111000,
    22'b0001111100001010001111,
    22'b0001110110100011110110,
    22'b0001101110101110000101,
    22'b0001101000010100011111,
    22'b0001100100011110101110,
    22'b0001011111110101110001,
    22'b0001011100011110101110,
    22'b0001011001011100001010,
    22'b0001010111000010100100,
    22'b0001010100001010001111,
    22'b0001001111000010100100,
    22'b0001001001110000101001,
    22'b0001000100010100011111,
    22'b0000111111101011100001,
    22'b0000111000111101011100,
    22'b0000110100000000000000,
    22'b0000101110100011110110,
    22'b0000101001010001111011,
    22'b0000100010111000010100,
    22'b0000011110101110000101,
    22'b0000011010111000010100,
    22'b0000011000011110101110,
    22'b0000010111001100110011,
    22'b0000010110100011110110,
    22'b0000010110000101001000,
    22'b0000010100010100011111,
    22'b0000010011100001010010,
    22'b0000010011110101110001,
    22'b0000010101000111101100,
    22'b0000010111110101110001,
    22'b0000011100000000000000,
    22'b0000100100110011001101,
    22'b0000101100011110101110,
    22'b0000110100110011001101,
    22'b0000111101011100001010,
    22'b0001000111101011100001,
    22'b0001001101100110011010,
    22'b0001010000010100011111,
    22'b0001010000000000000000,
    22'b0001001100010100011111,
    22'b0001001000010100011111,
    22'b0001000100101000111101,
    22'b0001000001010001111011,
    22'b0000111110100011110110,
    22'b0000111011110101110001,
    22'b0000111001110000101001,
    22'b0000110110111000010100,
    22'b0000110010101110000101,
    22'b0000101011001100110011,
    22'b0000100100001010001111,
    22'b0000011100001010001111,
    22'b0000010011110101110001,
    22'b0000001011110101110001,
    22'b0000000010000101001000,
    22'b1111111011100001010010,
    22'b1111110110001111010111,
    22'b1111110001110000101001,
    22'b1111101011100001010010,
    22'b1111100101011100001010,
    22'b1111011110100011110110,
    22'b1111010110100011110110,
    22'b1111001010111000010100,
    22'b1111000011001100110011,
    22'b1110111011001100110011,
    22'b1110110011001100110011,
    22'b1110101110011001100110,
    22'b1110101011000010100100,
    22'b1110101001011100001010,
    22'b1110101111000010100100,
    22'b1110110101111010111000,
    22'b1110111101111010111000,
    22'b1111000111110101110001,
    22'b1111010010000101001000,
    22'b1111011010011001100110,
    22'b1110111100011110101110,
    22'b1110110000000000000000,
    22'b1110101000101000111101,
    22'b1110100111001100110011,
    22'b1110100111000010100100,
    22'b1110100111010111000011,
    22'b1110100101110000101001,
    22'b1110100100010100011111,
    22'b1110101011100001010010,
    22'b1111000000101000111101,
    22'b1111001010101110000101,
    22'b1111001111010111000011,
    22'b1111010000101000111101,
    22'b1111001111101011100001,
    22'b1111001111000010100100,
    22'b1111001111001100110011,
    22'b1111001110000101001000,
    22'b1111001110001111010111,
    22'b1111001110111000010100,
    22'b1111001111001100110011,
    22'b1111001101111010111000,
    22'b1111001100001010001111,
    22'b1111001000010100011111,
    22'b1111000011100001010010,
    22'b1110111111001100110011,
    22'b1110111011000010100100,
    22'b1110110110000101001000,
    22'b1110110000111101011100,
    22'b1110101011100001010010,
    22'b1110100101100110011010,
    22'b1110011110001111010111,
    22'b1110010110101110000101,
    22'b1110001011010111000011,
    22'b1110000001011100001010,
    22'b1101111001000111101100,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101111000000000000000,
    22'b1110001000011110101110,
    22'b1110010111110101110001,
    22'b1110100101111010111000,
    22'b1110110001111010111000,
    22'b1110111101110000101001,
    22'b1111001010101110000101,
    22'b1111010001011100001010,
    22'b1111010011001100110011,
    22'b1111010001110000101001,
    22'b1111001110101110000101,
    22'b1111001000111101011100,
    22'b1111000011110101110001,
    22'b1110111110100011110110,
    22'b1110111000111101011100,
    22'b1110110001110000101001,
    22'b1110101100000000000000,
    22'b1110100101100110011010,
    22'b1110011110001111010111,
    22'b1110010101100110011010,
    22'b1110001000011110101110,
    22'b1101111101011100001010,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101111011001100110011,
    22'b1110000100011110101110,
    22'b1110001101010001111011,
    22'b1110010111110101110001,
    22'b1110011111000010100100,
    22'b1110100100011110101110,
    22'b1110101000101000111101,
    22'b1110101100001010001111,
    22'b1110101101110000101001,
    22'b1110101110001111010111,
    22'b1110101110000101001000,
    22'b1110101101011100001010,
    22'b1110101011101011100001,
    22'b1110101000110011001101,
    22'b1110100100110011001101,
    22'b1110100000010100011111,
    22'b1110011010011001100110,
    22'b1110010110011001100110,
    22'b1110010011010111000011,
    22'b1110010001010001111011,
    22'b1110010000111101011100,
    22'b1110010010111000010100,
    22'b1110010101111010111000,
    22'b1110011010001111010111,
    22'b1110011111000010100100,
    22'b1110100110001111010111,
    22'b1110101100011110101110,
    22'b1110110010111000010100,
    22'b1110111001110000101001,
    22'b1111000011001100110011,
    22'b1111001010100011110110,
    22'b1111010001111010111000,
    22'b1111011000101000111101,
    22'b1111100010000101001000,
    22'b1111101000111101011100,
    22'b1111101111101011100001,
    22'b1111110110000101001000,
    22'b1111111100000000000000,
    22'b0000000011101011100001,
    22'b0000001001000111101100,
    22'b0000001110101110000101,
    22'b0000010100010100011111,
    22'b0000011100001010001111,
    22'b0000100010001111010111,
    22'b0000101000010100011111,
    22'b0000101110111000010100,
    22'b0000110101100110011010,
    22'b0000111110001111010111,
    22'b0001000100010100011111,
    22'b0001001001111010111000,
    22'b0001001111001100110011,
    22'b0001010101100110011010,
    22'b0001011010000101001000,
    22'b0001011110111000010100,
    22'b0001100010111000010100,
    22'b0001100111010111000011,
    22'b0001101100011110101110,
    22'b0001101110000101001000,
    22'b0001101101111010111000,
    22'b0001101100001010001111,
    22'b0001101101011100001010,
    22'b0001101110000101001000,
    22'b0001101100010100011111,
    22'b0001101010111000010100,
    22'b0001101001000111101100,
    22'b0001100111100001010010,
    22'b0001100111110101110001,
    22'b0001100011010111000011,
    22'b0001100000001010001111,
    22'b0001011110111000010100,
    22'b0001100000001010001111,
    22'b0001100111100001010010,
    22'b0001101101111010111000,
    22'b0001101111110101110001,
    22'b0001110011001100110011,
    22'b0001111011010111000011,
    22'b0010000110011001100110,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010000111101011100001,
    22'b0001111101100110011010,
    22'b0001110000001010001111,
    22'b0001101001100110011010,
    22'b0001101001010001111011,
    22'b0001101111010111000011,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010000110000101001000,
    22'b0001011101100110011010,
    22'b0001001000011110101110,
    22'b0000111010111000010100,
    22'b0000101010000101001000,
    22'b0000101110011001100110,
    22'b0000101001011100001010,
    22'b0000011011001100110011,
    22'b1111111100110011001101,
    22'b1111111000010100011111,
    22'b1111111010001111010111,
    22'b0000000110000101001000,
    22'b0000001011100001010010,
    22'b1111111100010100011111,
    22'b1111011101111010111000,
    22'b1111000001100110011010,
    22'b1110110111000010100100,
    22'b1111010011000010100100,
    22'b1111001111110101110001,
    22'b1111001001100110011010,
    22'b1111001010101110000101,
    22'b1111010011010111000011,
    22'b1111011101110000101001,
    22'b1111101000010100011111,
    22'b1111110100101000111101,
    22'b1111111100010100011111,
    22'b0000000011010111000011,
    22'b0000000110011001100110,
    22'b1111111010001111010111,
    22'b1111101010101110000101,
    22'b1111011100101000111101,
    22'b1111010000101000111101,
    22'b1111000010101110000101,
    22'b1110110110111000010100,
    22'b1110100111000010100100,
    22'b1110010100111101011100,
    22'b1101111100001010001111,
    22'b1101110100010100011111,
    22'b1101111001100110011010,
    22'b1110110111001100110011,
    22'b1111101000110011001101,
    22'b1111101110100011110110,
    22'b1111101101100110011010,
    22'b1111110111100001010010,
    22'b1111111110000101001000,
    22'b1111111110100011110110,
    22'b1111111000001010001111,
    22'b1111110100001010001111,
    22'b1111110111101011100001,
    22'b1111110001011100001010,
    22'b1111100100000000000000,
    22'b1111001110001111010111,
    22'b1110111111010111000011,
    22'b1110110100011110101110,
    22'b1110110010011001100110,
    22'b1110101111100001010010,
    22'b1110110001100110011010,
    22'b1110111001011100001010,
    22'b1111000101010001111011,
    22'b1111010010011001100110,
    22'b1111010111010111000011,
    22'b1111010001010001111011,
    22'b1110111111110101110001,
    22'b1110110110111000010100,
    22'b1111000011101011100001,
    22'b1111001111010111000011,
    22'b1111010111010111000011,
    22'b1111011100010100011111,
    22'b1111011111000010100100,
    22'b1111100011000010100100,
    22'b1111100111101011100001,
    22'b1111101010100011110110,
    22'b1111101001111010111000,
    22'b1111101011110101110001,
    22'b1111110001100110011010,
    22'b1111110100000000000000,
    22'b0000000000001010001111,
    22'b0000000001111010111000,
    22'b0000000010111000010100,
    22'b0000000011001100110011,
    22'b0000000011001100110011,
    22'b0000000011000010100100,
    22'b0000000010100011110110,
    22'b0000000010011001100110,
    22'b0000000001111010111000,
    22'b0000000000110011001101,
    22'b1111111110100011110110,
    22'b1111111100101000111101,
    22'b1111111010111000010100,
    22'b1111111010000101001000,
    22'b1111111010000101001000,
    22'b1111111010011001100110,
    22'b1111111010100011110110,
    22'b1111111010001111010111,
    22'b1111111000111101011100,
    22'b1111110111100001010010,
    22'b1111110110001111010111,
    22'b1111110101100110011010,
    22'b1111110110000101001000,
    22'b1111110101111010111000,
    22'b1111110111110101110001,
    22'b1111111001111010111000,
    22'b1111111011101011100001,
    22'b1111111100110011001101,
    22'b1111111101110000101001,
    22'b1111111110011001100110,
    22'b1111111111100001010010,
    22'b0000000011010111000011,
    22'b0000000110011001100110,
    22'b0000001010100011110110,
    22'b0000001101000111101100,
    22'b0000001111010111000011,
    22'b0000010001011100001010,
    22'b0000010100011110101110,
    22'b0000010111001100110011,
    22'b0000011001111010111000,
    22'b0000011101110000101001,
    22'b0000011110000101001000,
    22'b0000100000000000000000,
    22'b0000100011100001010010,
    22'b0000100110100011110110,
    22'b0000101101000111101100,
    22'b0000110100011110101110,
    22'b0000111101111010111000,
    22'b0000111111001100110011,
    22'b0001001010000101001000,
    22'b0001010011001100110011,
    22'b0001010111100001010010,
    22'b0001011000001010001111,
    22'b0001011010101110000101,
    22'b0001011000000000000000,
    22'b0001010110111000010100,
    22'b0001011010000101001000,
    22'b0001011000010100011111,
    22'b0001011001010001111011,
    22'b0001011001100110011010,
    22'b0001011000101000111101,
    22'b0001010000010100011111,
    22'b0001001101110000101001,
    22'b0001001110101110000101,
    22'b0001001100111101011100,
    22'b0001001010111000010100,
    22'b0001001001100110011010,
    22'b0001001001011100001010,
    22'b0001001010000101001000,
    22'b0001001100110011001101,
    22'b0001010001000111101100,
    22'b0001010011001100110011,
    22'b0001010010011001100110,
    22'b0001010010001111010111,
    22'b0001010010011001100110,
    22'b0001010010011001100110,
    22'b0001010011001100110011,
    22'b0001010110011001100110,
    22'b0001011010001111010111,
    22'b0001011100001010001111,
    22'b0001011101000111101100,
    22'b0001011110111000010100,
    22'b0001100000011110101110,
    22'b0001100001010001111011,
    22'b0001100001100110011010,
    22'b0001100001100110011010,
    22'b0001100010001111010111,
    22'b0001100000110011001101,
    22'b0001011101110000101001,
    22'b0001011011110101110001,
    22'b0001011010011001100110,
    22'b0001011001100110011010,
    22'b0001011001000111101100,
    22'b0001011000101000111101,
    22'b0001010111101011100001,
    22'b0001010101100110011010,
    22'b0001010011001100110011,
    22'b0001010000101000111101,
    22'b0001001011100001010010,
    22'b0001000101111010111000,
    22'b0001001010111000010100,
    22'b0001001010000101001000,
    22'b0001000011010111000011,
    22'b0000111100101000111101,
    22'b0000110111101011100001,
    22'b0000110111101011100001,
    22'b0000110111001100110011,
    22'b0000110101110000101001,
    22'b0000110100011110101110,
    22'b0000110100011110101110,
    22'b0000110101110000101001,
    22'b0000110100011110101110,
    22'b0000110001010001111011,
    22'b0000101111101011100001,
    22'b0000110000000000000000,
    22'b0000110010011001100110,
    22'b0000110111110101110001,
    22'b0000111010100011110110,
    22'b0000110110101110000101,
    22'b0000110011010111000011,
    22'b0000110011010111000011,
    22'b0000110101111010111000,
    22'b0000110110001111010111,
    22'b0000110011001100110011,
    22'b0000101101010001111011,
    22'b0000100111101011100001,
    22'b0000011110000101001000,
    22'b0000010010111000010100,
    22'b0000010001011100001010,
    22'b0000001011001100110011,
    22'b0000001011110101110001,
    22'b0000010000001010001111,
    22'b0000010101100110011010,
    22'b0000010101010001111011,
    22'b0000010010011001100110,
    22'b0000010001000111101100,
    22'b0000010001110000101001,
    22'b0000010011100001010010,
    22'b0000010100101000111101,
    22'b0000010101110000101001,
    22'b0000010110001111010111,
    22'b0000010110100011110110,
    22'b0000010111010111000011,
    22'b0000011000011110101110,
    22'b0000011001011100001010,
    22'b0000011000101000111101,
    22'b0000010101110000101001,
    22'b0000010100011110101110,
    22'b0000010010000101001000,
    22'b0000001100001010001111,
    22'b0000000000101000111101,
    22'b1111110011110101110001,
    22'b1111101010101110000101,
    22'b1111100111100001010010,
    22'b1111101010011001100110,
    22'b1111110000101000111101,
    22'b1111110111100001010010,
    22'b1111111101000111101100,
    22'b0000000001100110011010,
    22'b0000000010011001100110,
    22'b0000000011100001010010,
    22'b0000000000111101011100,
    22'b1111111101011100001010,
    22'b1111111001100110011010,
    22'b1111110110011001100110,
    22'b1111110100101000111101,
    22'b1111110101000111101100,
    22'b1111110101010001111011,
    22'b1111110101010001111011,
    22'b1111110101010001111011,
    22'b1111110101110000101001,
    22'b1111110110000101001000,
    22'b1111110101111010111000,
    22'b1111110100110011001101,
    22'b1111110111100001010010,
    22'b1111110111010111000011,
    22'b1111110110111000010100,
    22'b1111110011100001010010,
    22'b1111110001110000101001,
    22'b1111110010011001100110,
    22'b1111100011110101110001,
    22'b1111011010000101001000,
    22'b1111011001110000101001,
    22'b1111010101110000101001,
    22'b1111010111100001010010,
    22'b1111011101111010111000,
    22'b1111100100110011001101,
    22'b1111101110001111010111,
    22'b1111111001110000101001,
    22'b1111111111000010100100,
    22'b0000000011101011100001,
    22'b0000000011110101110001,
    22'b0000000010100011110110,
    22'b0000000001111010111000,
    22'b0000000010100011110110,
    22'b0000000101100110011010,
    22'b0000001001111010111000,
    22'b0000001110100011110110,
    22'b0000010010000101001000,
    22'b0000010100101000111101,
    22'b0000010101100110011010,
    22'b0000010110000101001000,
    22'b0000011000011110101110,
    22'b0000100110001111010111,
    22'b0000101111001100110011,
    22'b0000110000011110101110,
    22'b0000101011010111000011,
    22'b0000100001010001111011,
    22'b0000011100010100011111,
    22'b0000011001100110011010,
    22'b0000011001010001111011,
    22'b0000100010101110000101,
    22'b0000101100111101011100,
    22'b0000100000001010001111,
    22'b0000001101100110011010,
    22'b0000001011001100110011,
    22'b0000010000000000000000,
    22'b0000010100010100011111,
    22'b0000011001111010111000,
    22'b0000011111001100110011,
    22'b0000100000001010001111,
    22'b0000011111010111000011,
    22'b0000011101010001111011,
    22'b0000011010000101001000,
    22'b0000011001100110011010,
    22'b0000011001011100001010,
    22'b0000011010000101001000,
    22'b0000100000000000000000,
    22'b0000100010100011110110,
    22'b0000011110001111010111,
    22'b0000011000110011001101,
    22'b0000010110111000010100,
    22'b0000010111101011100001,
    22'b0000010111110101110001,
    22'b0000010111000010100100,
    22'b0000010101000111101100,
    22'b0000010100000000000000,
    22'b0000010010111000010100,
    22'b0000010001111010111000,
    22'b0000010000110011001101,
    22'b0000001110111000010100,
    22'b0000001101010001111011,
    22'b0000001011101011100001,
    22'b0000001010011001100110,
    22'b0000001000111101011100,
    22'b0000001000001010001111,
    22'b0000000111100001010010,
    22'b0000000111000010100100,
    22'b0000000110100011110110,
    22'b0000000110001111010111,
    22'b0000000101111010111000,
    22'b0000000101111010111000,
    22'b0000000101011100001010,
    22'b0000000100101000111101,
    22'b0000000100000000000000,
    22'b0000000011100001010010,
    22'b0000000011010111000011,
    22'b0000000011110101110001,
    22'b0000000100010100011111,
    22'b0000000101000111101100,
    22'b0000000110011001100110,
    22'b0000000111110101110001,
    22'b0000001000110011001101,
    22'b0000001001110000101001,
    22'b0000001010011001100110,
    22'b0000001011001100110011,
    22'b0000001100001010001111,
    22'b0000001100111101011100,
    22'b0000001101100110011010,
    22'b0000001110000101001000,
    22'b0000001110100011110110,
    22'b0000001110100011110110,
    22'b0000001100011110101110,
    22'b0000000111110101110001,
    22'b0000001000001010001111,
    22'b0000000101110000101001,
    22'b0000000100000000000000,
    22'b0000000010100011110110,
    22'b0000000010011001100110,
    22'b0000000010101110000101,
    22'b0000000011010111000011,
    22'b0000000100010100011111,
    22'b0000000100110011001101,
    22'b0000000100111101011100,
    22'b0000000100111101011100,
    22'b0000000100110011001101,
    22'b0000000100101000111101,
    22'b0000000100011110101110,
    22'b0000000100000000000000,
    22'b0000000100001010001111,
    22'b0000000100110011001101,
    22'b0000000110001111010111,
    22'b0000001000000000000000,
    22'b0000001000101000111101,
    22'b0000001001010001111011,
    22'b0000001010001111010111,
    22'b0000001011001100110011,
    22'b0000001011110101110001,
    22'b0000001011110101110001,
    22'b0000001011001100110011,
    22'b0000001000110011001101,
    22'b0000000111001100110011,
    22'b0000000111001100110011,
    22'b0000000111001100110011,
    22'b0000000110001111010111,
    22'b0000000100101000111101,
    22'b0000000010101110000101,
    22'b0000000001010001111011,
    22'b1111111111101011100001,
    22'b1111111110001111010111,
    22'b1111111101010001111011,
    22'b1111111100110011001101,
    22'b1111111100000000000000,
    22'b1111111010011001100110,
    22'b1111111001110000101001,
    22'b1111111001100110011010,
    22'b1111111001100110011010,
    22'b1111111001011100001010,
    22'b1111111001000111101100,
    22'b1111111000011110101110,
    22'b1111110111001100110011,
    22'b1111110101100110011010,
    22'b1111110011100001010010,
    22'b1111110010001111010111,
    22'b1111110001010001111011,
    22'b1111110000011110101110,
    22'b1111101110111000010100,
    22'b1111101101011100001010,
    22'b1111101011101011100001,
    22'b1111101001110000101001,
    22'b1111100111001100110011,
    22'b1111100101010001111011,
    22'b1111100011101011100001,
    22'b1111100010100011110110,
    22'b1111100001110000101001,
    22'b1111100000101000111101,
    22'b1111011111001100110011,
    22'b1111011101100110011010,
    22'b1111011100011110101110,
    22'b1111011011100001010010,
    22'b1111011010101110000101,
    22'b1111011010000101001000,
    22'b1111011010000101001000,
    22'b1111011010001111010111,
    22'b1111011010011001100110,
    22'b1111011010001111010111,
    22'b1111011001100110011010,
    22'b1111011001000111101100,
    22'b1111010111110101110001,
    22'b1111010110100011110110,
    22'b1111010101011100001010,
    22'b1111010100000000000000,
    22'b1111010010011001100110,
    22'b1111010000110011001101,
    22'b1111010000011110101110,
    22'b1111010000101000111101,
    22'b1111001111010111000011,
    22'b1111001001011100001010,
    22'b1111001000111101011100,
    22'b1111001001011100001010,
    22'b1111001011001100110011,
    22'b1111001101111010111000,
    22'b1111001110111000010100,
    22'b1111010000001010001111,
    22'b1111010010000101001000,
    22'b1111010100011110101110,
    22'b1111011100000000000000,
    22'b1111011111001100110011,
    22'b1111100001000111101100,
    22'b1111100010100011110110,
    22'b1111100011110101110001,
    22'b1111100101010001111011,
    22'b1111100110001111010111,
    22'b1111100110101110000101,
    22'b1111100111010111000011,
    22'b1111101000001010001111,
    22'b1111101000110011001101,
    22'b1111101001100110011010,
    22'b1111101010101110000101,
    22'b1111101100001010001111,
    22'b1111101111001100110011,
    22'b1111110101110000101001,
    22'b0000001000011110101110,
    22'b0000001111010111000011,
    22'b0000010000001010001111,
    22'b0000000001011100001010,
    22'b1111111110101110000101,
    22'b0000000010111000010100,
    22'b0000000111101011100001,
    22'b0000000110100011110110,
    22'b1111111010000101001000,
    22'b1111110011101011100001,
    22'b1111110000111101011100,
    22'b1111110010101110000101,
    22'b1111111010000101001000,
    22'b1111110111001100110011,
    22'b1111110010101110000101,
    22'b1111101110101110000101,
    22'b1111101011001100110011,
    22'b1111100111010111000011,
    22'b1111100110000101001000,
    22'b1111100101010001111011,
    22'b1111100101000111101100,
    22'b1111100101010001111011,
    22'b1111100101011100001010,
    22'b1111100101110000101001,
    22'b1111100110100011110110,
    22'b1111101000000000000000,
    22'b1111101001100110011010,
    22'b1111101011101011100001,
    22'b1111101110100011110110,
    22'b1111110000110011001101,
    22'b1111101110111000010100,
    22'b1111101101110000101001,
    22'b1111110011010111000011,
    22'b1111111110000101001000,
    22'b0000000101000111101100,
    22'b0000010110011001100110,
    22'b0000001110100011110110,
    22'b0000001000110011001101,
    22'b0000000110100011110110,
    22'b0000001011000010100100,
    22'b0000010001000111101100,
    22'b0000011111100001010010,
    22'b0000110001100110011010,
    22'b0001000011000010100100,
    22'b0001010100101000111101,
    22'b0001011101110000101001,
    22'b0001011110011001100110,
    22'b0001011100011110101110,
    22'b0001010001011100001010,
    22'b0001000000011110101110,
    22'b0000101010111000010100,
    22'b0000011100010100011111,
    22'b0000010000010100011111,
    22'b0000001000101000111101,
    22'b0000000101010001111011,
    22'b0000000100010100011111,
    22'b0000000100010100011111,
    22'b0000000100010100011111,
    22'b0000000011110101110001,
    22'b0000000010111000010100,
    22'b0000000000110011001101,
    22'b1111111110101110000101,
    22'b1111111100110011001101,
    22'b1111111011001100110011,
    22'b1111111010000101001000,
    22'b1111111001010001111011,
    22'b1111111001000111101100,
    22'b1111111000111101011100,
    22'b1111111000011110101110,
    22'b1111110111100001010010,
    22'b1111110101111010111000,
    22'b1111110100011110101110,
    22'b1111110011010111000011,
    22'b1111110010100011110110,
    22'b1111110001011100001010,
    22'b1111101111110101110001,
    22'b1111101110011001100110,
    22'b1111101100010100011111,
    22'b1111101001011100001010,
    22'b1111100101100110011010,
    22'b1111100010101110000101,
    22'b1111011111101011100001,
    22'b1111011100101000111101,
    22'b1111011001110000101001,
    22'b1111010111010111000011,
    22'b1111010111000010100100,
    22'b1111011000011110101110,
    22'b1111011011010111000011,
    22'b1111100000111101011100,
    22'b1111100101100110011010,
    22'b1111101010001111010111,
    22'b1111101110011001100110,
    22'b1111110001111010111000,
    22'b1111110110001111010111,
    22'b1111111001011100001010,
    22'b1111111101110000101001,
    22'b0000000011000010100100,
    22'b0000001110000101001000,
    22'b0000010111101011100001,
    22'b0000100000011110101110,
    22'b0000100111110101110001,
    22'b0000101111010111000011,
    22'b0000110110111000010100,
    22'b0000111001011100001010,
    22'b0000111100011110101110,
    22'b0000111101011100001010,
    22'b0000111100000000000000,
    22'b0000111011000010100100,
    22'b0000110111100001010010,
    22'b0000110100011110101110,
    22'b0000110001000111101100,
    22'b0000101101010001111011,
    22'b0000101001110000101001,
    22'b0000100101111010111000,
    22'b0000100100000000000000,
    22'b0000100010100011110110,
    22'b0000100001110000101001,
    22'b0000100001000111101100,
    22'b0000100001010001111011,
    22'b0000100001000111101100,
    22'b0000100000101000111101,
    22'b0000011111100001010010,
    22'b0000011100110011001101,
    22'b0000011010001111010111,
    22'b0000010111100001010010,
    22'b0000010100111101011100,
    22'b0000010010101110000101,
    22'b0000010000000000000000,
    22'b0000001110011001100110,
    22'b0000001100101000111101,
    22'b0000001001110000101001,
    22'b0000000111001100110011,
    22'b0000000100010100011111,
    22'b0000000011001100110011,
    22'b0000000010111000010100,
    22'b0000000011100001010010,
    22'b0000000101000111101100,
    22'b0000000111001100110011,
    22'b0000001000010100011111,
    22'b0000001000101000111101,
    22'b0000001000101000111101,
    22'b0000001000001010001111,
    22'b0000000111000010100100,
    22'b0000000110011001100110,
    22'b0000000110000101001000,
    22'b0000000101111010111000,
    22'b0000000110000101001000,
    22'b0000000110100011110110,
    22'b0000000110101110000101,
    22'b0000000110100011110110,
    22'b0000000110011001100110,
    22'b0000000101111010111000,
    22'b0000000011110101110001,
    22'b0000000100101000111101,
    22'b0000000100110011001101,
    22'b0000000100001010001111,
    22'b0000000110000101001000,
    22'b0000000110100011110110,
    22'b0000000111001100110011,
    22'b0000001000001010001111,
    22'b0000001000101000111101,
    22'b0000001001000111101100,
    22'b0000001000110011001101,
    22'b0000000111110101110001,
    22'b0000000111001100110011,
    22'b0000000110100011110110,
    22'b0000000101010001111011,
    22'b0000000001111010111000,
    22'b1111111101110000101001,
    22'b1111111110100011110110,
    22'b1111111111101011100001,
    22'b0000000000111101011100,
    22'b0000000001010001111011,
    22'b0000000001010001111011,
    22'b0000000000101000111101,
    22'b0000000000010100011111,
    22'b0000000000000000000000,
    22'b0000000000011110101110,
    22'b0000000001111010111000,
    22'b0000000101000111101100,
    22'b0000000111110101110001,
    22'b0000001010101110000101,
    22'b0000001110001111010111,
    22'b0000010011010111000011,
    22'b0000010110101110000101,
    22'b0000011001111010111000,
    22'b0000011111101011100001,
    22'b0000101010011001100110,
    22'b0000110001000111101100,
    22'b0000110101000111101100,
    22'b0000111001100110011010,
    22'b0000111101010001111011,
    22'b0001000000000000000000,
    22'b0001000001011100001010,
    22'b0001000010001111010111,
    22'b0001000001010001111011,
    22'b0000111111000010100100,
    22'b0000111011110101110001,
    22'b0000111100011110101110,
    22'b0000111100010100011111,
    22'b0000111000001010001111,
    22'b0000110111010111000011,
    22'b0000110010101110000101,
    22'b0000110000111101011100,
    22'b0000110000110011001101,
    22'b0000100100110011001101,
    22'b0000010101000111101100,
    22'b0000000011101011100001,
    22'b1111110001110000101001,
    22'b1111100000000000000000,
    22'b1111001010100011110110,
    22'b1110111100110011001101,
    22'b1110110000001010001111,
    22'b1110100101100110011010,
    22'b1110011011100001010010,
    22'b1110010101011100001010,
    22'b1110001111110101110001,
    22'b1110001011010111000011,
    22'b1110001010000101001000,
    22'b1110001110000101001000,
    22'b1110010010111000010100,
    22'b1110010111100001010010,
    22'b1110100000001010001111,
    22'b1110100111110101110001,
    22'b1110101110101110000101,
    22'b1110110100101000111101,
    22'b1110111001110000101001,
    22'b1111000000000000000000,
    22'b1111000100001010001111,
    22'b1111001000001010001111,
    22'b1111001011100001010010,
    22'b1111001111010111000011,
    22'b1111010010000101001000,
    22'b1111010101100110011010,
    22'b1111011010100011110110,
    22'b1111100000110011001101,
    22'b1111101010100011110110,
    22'b1111110010001111010111,
    22'b1111111010001111010111,
    22'b0000000010100011110110,
    22'b0000001110001111010111,
    22'b0000010111000010100100,
    22'b0000011111100001010010,
    22'b0000101000000000000000,
    22'b0000110000101000111101,
    22'b0000111011000010100100,
    22'b0001000001110000101001,
    22'b0001000111001100110011,
    22'b0001001100001010001111,
    22'b0001010001011100001010,
    22'b0001011001000111101100,
    22'b0001011111010111000011,
    22'b0001100101011100001010,
    22'b0001100110101110000101,
    22'b0001011101010001111011,
    22'b0001000011110101110001,
    22'b0000110000010100011111,
    22'b0000100000110011001101,
    22'b0000010101010001111011,
    22'b0000001101010001111011,
    22'b0000000111100001010010,
    22'b0000000111100001010010,
    22'b0000001100110011001101,
    22'b0000010111100001010010,
    22'b0000101100111101011100,
    22'b0001000000110011001101,
    22'b0001010110011001100110,
    22'b0001101101000111101100,
    22'b0010000100001010001111,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0001101101000111101100,
    22'b0001010010000101001000,
    22'b0001001000010100011111,
    22'b0001000011001100110011,
    22'b0001000001110000101001,
    22'b0001000100001010001111,
    22'b0001000101110000101001,
    22'b0001001001110000101001,
    22'b0001001111110101110001,
    22'b0001010111110101110001,
    22'b0001100010011001100110,
    22'b0001100110001111010111,
    22'b0001101001111010111000,
    22'b0001101101110000101001,
    22'b0001101110011001100110,
    22'b0001101100011110101110,
    22'b0001101011000010100100,
    22'b0001101101100110011010,
    22'b0001101110100011110110,
    22'b0001101100110011001101,
    22'b0001101000010100011111,
    22'b0001100100010100011111,
    22'b0001100001111010111000,
    22'b0001011111101011100001,
    22'b0001011011110101110001,
    22'b0001011000110011001101,
    22'b0001010101110000101001,
    22'b0001010010001111010111,
    22'b0001001101011100001010,
    22'b0001000110011001100110,
    22'b0001000010011001100110,
    22'b0000111111101011100001,
    22'b0000111100111101011100,
    22'b0000111001110000101001,
    22'b0000111000000000000000,
    22'b0000110110001111010111,
    22'b0000110100011110101110,
    22'b0000110001011100001010,
    22'b0000101101110000101001,
    22'b0000101101010001111011,
    22'b0000101100111101011100,
    22'b0000101011000010100100,
    22'b0000101000000000000000,
    22'b0000100100001010001111,
    22'b0000100010000101001000,
    22'b0000011111100001010010,
    22'b0000011100110011001101,
    22'b0000011011001100110011,
    22'b0000011001000111101100,
    22'b0000010110001111010111,
    22'b0000001111101011100001,
    22'b0000001000011110101110,
    22'b1111111111010111000011,
    22'b1111110011110101110001,
    22'b1111100000000000000000,
    22'b1111001101100110011010,
    22'b1110111001011100001010,
    22'b1110100101011100001010,
    22'b1110001110011001100110,
    22'b1110000001010001111011,
    22'b1101111000001010001111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101111000011110101110,
    22'b1101111011101011100001,
    22'b1101111101000111101100,
    22'b1110000110001111010111,
    22'b1110010001010001111011,
    22'b1110010110011001100110,
    22'b1110011111001100110011,
    22'b1110100000101000111101,
    22'b1110011110111000010100,
    22'b1110011001111010111000,
    22'b1110001110111000010100,
    22'b1110000111001100110011,
    22'b1110000001000111101100,
    22'b1101110111010111000011,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1110000111000010100100,
    22'b1110100111000010100100,
    22'b1110111000000000000000,
    22'b1111000000101000111101,
    22'b1111000100110011001101,
    22'b1111001001011100001010,
    22'b1111001101000111101100,
    22'b1111010001000111101100,
    22'b1111010100010100011111,
    22'b1111010111100001010010,
    22'b1111011010011001100110,
    22'b1111011110001111010111,
    22'b1111011111100001010010,
    22'b1111011101010001111011,
    22'b1111011010100011110110,
    22'b1111011100111101011100,
    22'b1111011111101011100001,
    22'b1111100010001111010111,
    22'b1111100101100110011010,
    22'b1111101000000000000000,
    22'b1111101010000101001000,
    22'b1111101100000000000000,
    22'b1111101110001111010111,
    22'b1111101111110101110001,
    22'b1111110001000111101100,
    22'b1111110010000101001000,
    22'b1111110010101110000101,
    22'b1111110011001100110011,
    22'b1111110011000010100100,
    22'b1111110011101011100001,
    22'b1111110100010100011111,
    22'b1111110100001010001111,
    22'b1111110001100110011010,
    22'b1111101100000000000000,
    22'b1111101001000111101100,
    22'b1111100110011001100110,
    22'b1111100011000010100100,
    22'b1111011110000101001000,
    22'b1111011000010100011111,
    22'b1111010000000000000000,
    22'b1111000100000000000000,
    22'b1110111010101110000101,
    22'b1110110011101011100001,
    22'b1110110000111101011100,
    22'b1110101110100011110110,
    22'b1110111010101110000101,
    22'b1111001011010111000011,
    22'b1111010101100110011010,
    22'b1111011100011110101110,
    22'b1111100101110000101001,
    22'b1111101011000010100100,
    22'b1111101111001100110011,
    22'b1111110010100011110110,
    22'b1111110011110101110001,
    22'b1111110100101000111101,
    22'b1111110100011110101110,
    22'b1111110010101110000101,
    22'b1111110000110011001101,
    22'b1111101111001100110011,
    22'b1111101101110000101001,
    22'b1111101100110011001101,
    22'b1111101100001010001111,
    22'b1111101011000010100100,
    22'b1111101010000101001000,
    22'b1111101000101000111101,
    22'b1111100111101011100001,
    22'b1111100111010111000011,
    22'b1111101001000111101100,
    22'b1111101010100011110110,
    22'b1111101011110101110001,
    22'b1111101101100110011010,
    22'b1111101111100001010010,
    22'b1111110000111101011100,
    22'b1111110010100011110110,
    22'b1111110011100001010010,
    22'b1111110101000111101100,
    22'b1111110110100011110110,
    22'b1111110111001100110011,
    22'b1111110111101011100001,
    22'b1111111000110011001101,
    22'b1111111100111101011100,
    22'b1111111110001111010111,
    22'b0000000000001010001111,
    22'b0000000001110000101001,
    22'b0000000011010111000011,
    22'b0000000100101000111101,
    22'b0000000110001111010111,
    22'b0000000111000010100100,
    22'b0000000111110101110001,
    22'b0000001000101000111101,
    22'b0000001001011100001010,
    22'b0000001001111010111000,
    22'b0000001010011001100110,
    22'b0000001010111000010100,
    22'b0000001011000010100100,
    22'b0000001011100001010010,
    22'b0000001011110101110001,
    22'b0000001100001010001111,
    22'b0000001100101000111101,
    22'b0000001101000111101100,
    22'b0000001101100110011010,
    22'b0000001101111010111000,
    22'b0000001110001111010111,
    22'b0000001110100011110110,
    22'b0000001110111000010100,
    22'b0000001111010111000011,
    22'b0000001111110101110001,
    22'b0000010000001010001111,
    22'b0000010000011110101110,
    22'b0000010000110011001101,
    22'b0000010001011100001010,
    22'b0000010001100110011010,
    22'b0000010001110000101001,
    22'b0000010001100110011010,
    22'b0000010001110000101001,
    22'b0000010010001111010111,
    22'b0000010010100011110110,
    22'b0000010010101110000101,
    22'b0000010010011001100110,
    22'b0000010001111010111000,
    22'b0000010001011100001010,
    22'b0000010001000111101100,
    22'b0000010000101000111101,
    22'b0000010000010100011111,
    22'b0000001111101011100001,
    22'b0000001111001100110011,
    22'b0000001110011001100110,
    22'b0000001110000101001000,
    22'b0000001101111010111000,
    22'b0000001101110000101001,
    22'b0000001101110000101001,
    22'b0000001101110000101001,
    22'b0000001101110000101001,
    22'b0000001101111010111000,
    22'b0000001101111010111000,
    22'b0000001101110000101001,
    22'b0000001101100110011010,
    22'b0000001101000111101100,
    22'b0000001100110011001101,
    22'b0000001100011110101110,
    22'b0000001100001010001111,
    22'b0000001011101011100001,
    22'b0000001011100001010010,
    22'b0000001011010111000011,
    22'b0000001011010111000011,
    22'b0000001011001100110011,
    22'b0000001011001100110011,
    22'b0000001011001100110011,
    22'b0000001011000010100100,
    22'b0000001010111000010100,
    22'b0000001010101110000101,
    22'b0000001010100011110110,
    22'b0000001010011001100110,
    22'b0000001010000101001000,
    22'b0000001000010100011111,
    22'b0000000011101011100001,
    22'b1111111111100001010010,
    22'b1111111110011001100110,
    22'b1111111101110000101001,
    22'b1111111100111101011100,
    22'b1111111011110101110001,
    22'b1111111011110101110001,
    22'b1111111100000000000000,
    22'b1111111100000000000000,
    22'b1111111011110101110001,
    22'b1111111011010111000011,
    22'b1111111010100011110110,
    22'b1111111001010001111011,
    22'b1111110111010111000011,
    22'b1111110101110000101001,
    22'b1111110100011110101110,
    22'b1111110011100001010010,
    22'b1111110001110000101001,
    22'b1111101111000010100100,
    22'b1111101101000111101100,
    22'b1111101100010100011111,
    22'b1111101011000010100100,
    22'b1111101010001111010111,
    22'b1111101010000101001000,
    22'b1111101001000111101100,
    22'b1111101000011110101110,
    22'b1111100111101011100001,
    22'b1111101000010100011111,
    22'b1111101010100011110110,
    22'b1111101101110000101001,
    22'b1111110000101000111101,
    22'b1111110011001100110011,
    22'b0000000000001010001111,
    22'b0000000010101110000101,
    22'b0000001100010100011111,
    22'b0000011101010001111011,
    22'b0000110100110011001101,
    22'b0000111110100011110110,
    22'b0000110010011001100110,
    22'b0000101111000010100100,
    22'b0000110011001100110011,
    22'b0000111001111010111000,
    22'b0001000001011100001010,
    22'b0001000000110011001101,
    22'b0000111010000101001000,
    22'b0000110001010001111011,
    22'b0000101100000000000000,
    22'b0000101100001010001111,
    22'b0000101101011100001010,
    22'b0000101101011100001010,
    22'b0000101011000010100100,
    22'b0000101001110000101001,
    22'b0000101000110011001101,
    22'b0000100111001100110011,
    22'b0000100110000101001000,
    22'b0000100101100110011010,
    22'b0000100100011110101110,
    22'b0000100011010111000011,
    22'b0000100010011001100110,
    22'b0000100001010001111011,
    22'b0000011111110101110001,
    22'b0000011100110011001101,
    22'b0000001001110000101001,
    22'b1111011001000111101100,
    22'b1110101001100110011010,
    22'b1110011110011001100110,
    22'b1110110011000010100100,
    22'b1111000110011001100110,
    22'b1111010110100011110110,
    22'b1111100010001111010111,
    22'b1111101111001100110011,
    22'b1111111000000000000000,
    22'b1111111100010100011111,
    22'b1111111011100001010010,
    22'b1111110110011001100110,
    22'b1111110011110101110001,
    22'b1111110011110101110001,
    22'b1111110011100001010010,
    22'b1111110011110101110001,
    22'b1111110110000101001000,
    22'b1111110111110101110001,
    22'b1111111001010001111011,
    22'b1111111010001111010111,
    22'b1111111010000101001000,
    22'b1111111010000101001000,
    22'b1111111010001111010111,
    22'b1111111000000000000000,
    22'b1111111001111010111000,
    22'b1111111010111000010100,
    22'b1111111011101011100001,
    22'b1111111100101000111101,
    22'b1111111101110000101001,
    22'b0000000000000000000000,
    22'b0000000010101110000101,
    22'b0000000110000101001000,
    22'b0000001000110011001101,
    22'b0000001011110101110001,
    22'b0000001110001111010111,
    22'b0000001111101011100001,
    22'b0000010001100110011010,
    22'b0000010011000010100100,
    22'b0000010010001111010111,
    22'b0000001110011001100110,
    22'b0000001011001100110011,
    22'b0000000011100001010010,
    22'b1111110010000101001000,
    22'b1111101101111010111000,
    22'b1111110110101110000101,
    22'b1111110111110101110001,
    22'b1111110100111101011100,
    22'b1111110001111010111000,
    22'b1111110010101110000101,
    22'b1111110010011001100110,
    22'b1111110001010001111011,
    22'b1111110000111101011100,
    22'b1111110000110011001101,
    22'b1111110000010100011111,
    22'b1111101111110101110001,
    22'b1111101111001100110011,
    22'b1111101110111000010100,
    22'b1111101111000010100100,
    22'b1111110000101000111101,
    22'b1111110010101110000101,
    22'b1111110100000000000000,
    22'b1111110101010001111011,
    22'b1111110101110000101001,
    22'b1111110110000101001000,
    22'b1111110110100011110110,
    22'b1111110110111000010100,
    22'b1111110110101110000101,
    22'b1111110110011001100110,
    22'b1111110110000101001000,
    22'b1111110101010001111011,
    22'b1111110100110011001101,
    22'b1111110100010100011111,
    22'b1111110011101011100001,
    22'b1111110011000010100100,
    22'b1111110010101110000101,
    22'b1111110011000010100100,
    22'b1111110101000111101100,
    22'b1111110100101000111101,
    22'b1111110010011001100110,
    22'b1111101111101011100001,
    22'b1111101111000010100100,
    22'b1111101111110101110001,
    22'b1111110000101000111101,
    22'b1111110001000111101100,
    22'b1111110000110011001101,
    22'b1111101111010111000011,
    22'b1111101110111000010100,
    22'b1111110000010100011111,
    22'b1111110000011110101110,
    22'b1111110000001010001111,
    22'b1111101110111000010100,
    22'b1111101110100011110110,
    22'b1111101101000111101100,
    22'b1111101010011001100110,
    22'b1111101000010100011111,
    22'b1111101001111010111000,
    22'b1111101001111010111000,
    22'b1111100111101011100001,
    22'b1111100101110000101001,
    22'b1111100101111010111000,
    22'b1111100111110101110001,
    22'b1111100111110101110001,
    22'b1111101000001010001111,
    22'b1111101000010100011111,
    22'b1111101000111101011100,
    22'b1111101000000000000000,
    22'b1111100111000010100100,
    22'b1111100110001111010111,
    22'b1111100100001010001111,
    22'b1111100010000101001000,
    22'b1111011111101011100001,
    22'b1111011001110000101001,
    22'b1111011000101000111101,
    22'b1111100001011100001010,
    22'b1111110010001111010111,
    22'b0000000010000101001000,
    22'b0000000100110011001101,
    22'b0000000010101110000101,
    22'b1111111111110101110001,
    22'b1111111001100110011010,
    22'b1111111011101011100001,
    22'b1111111011100001010010,
    22'b1111111000110011001101,
    22'b1111111011000010100100,
    22'b1111111111001100110011,
    22'b0000000010111000010100,
    22'b0000000110101110000101,
    22'b0000001010111000010100,
    22'b0000010000001010001111,
    22'b0000010011010111000011,
    22'b0000010101000111101100,
    22'b0000010110100011110110,
    22'b0000010110111000010100,
    22'b0000010110000101001000,
    22'b0000010101100110011010,
    22'b0000010100101000111101,
    22'b0000010001110000101001,
    22'b0000001110011001100110,
    22'b0000001100001010001111,
    22'b0000001010011001100110,
    22'b0000000111010111000011,
    22'b0000001000110011001101,
    22'b0000010000010100011111,
    22'b0000010001011100001010,
    22'b0000010000000000000000,
    22'b0000010011101011100001,
    22'b0000011011100001010010,
    22'b0000100011100001010010,
    22'b0000100010111000010100,
    22'b0000100001011100001010,
    22'b0000100010111000010100,
    22'b0000100101100110011010,
    22'b0000101011101011100001,
    22'b0000100111100001010010,
    22'b0000100101010001111011,
    22'b0000100001110000101001,
    22'b0000011111110101110001,
    22'b0000011011100001010010,
    22'b0000010011000010100100,
    22'b0000001011001100110011,
    22'b0000000011001100110011,
    22'b1111111100110011001101,
    22'b1111111110100011110110,
    22'b0000000010011001100110,
    22'b0000000100000000000000,
    22'b0000000110100011110110,
    22'b0000001100010100011111,
    22'b0000001111001100110011,
    22'b0000001111101011100001,
    22'b0000001110100011110110,
    22'b0000001100010100011111,
    22'b0000001001111010111000,
    22'b0000000101000111101100,
    22'b1111111110000101001000,
    22'b1111110011000010100100,
    22'b1111100111110101110001,
    22'b1111100010001111010111,
    22'b1111100100111101011100,
    22'b1111101010111000010100,
    22'b1111110000000000000000,
    22'b1111110100010100011111,
    22'b1111111000001010001111,
    22'b1111111000011110101110,
    22'b1111110001100110011010,
    22'b1111101110100011110110,
    22'b1111101100001010001111,
    22'b1111101011000010100100,
    22'b1111101100000000000000,
    22'b1111110010100011110110,
    22'b1111000110111000010100,
    22'b1110110001111010111000,
    22'b1110101001110000101001,
    22'b1110100111010111000011,
    22'b1110101110001111010111,
    22'b1110111000011110101110,
    22'b1111001110011001100110,
    22'b1111011000110011001101,
    22'b1111011101000111101100,
    22'b1111100001111010111000,
    22'b1111100000001010001111,
    22'b1111011110111000010100,
    22'b1111100100000000000000,
    22'b1111101010100011110110,
    22'b1111101010100011110110,
    22'b1111100011110101110001,
    22'b1111100000010100011111,
    22'b1111011111101011100001,
    22'b1111100010001111010111,
    22'b1111100101011100001010,
    22'b1111100110101110000101,
    22'b1111100111101011100001,
    22'b1111101000011110101110,
    22'b1111101001111010111000,
    22'b1111101111000010100100,
    22'b1111110011001100110011,
    22'b1111110101000111101100,
    22'b1111110101111010111000,
    22'b1111110111100001010010,
    22'b1111111000101000111101,
    22'b1111111001110000101001,
    22'b1111111010100011110110,
    22'b1111111011101011100001,
    22'b1111111101010001111011,
    22'b1111111111000010100100,
    22'b0000000001000111101100,
    22'b0000000011001100110011,
    22'b0000000101010001111011,
    22'b0000001000111101011100,
    22'b0000001100011110101110,
    22'b0000001111101011100001,
    22'b0000010011100001010010,
    22'b0000011000110011001101,
    22'b0000100000001010001111,
    22'b0000100101010001111011,
    22'b0000101100000000000000,
    22'b0000110001100110011010,
    22'b0000110100110011001101,
    22'b0000110100101000111101,
    22'b0000110011001100110011,
    22'b0000110000111101011100,
    22'b0000101110000101001000,
    22'b0000101010100011110110,
    22'b0000100101110000101001,
    22'b0000100001100110011010,
    22'b0000011100101000111101,
    22'b0000010110100011110110,
    22'b0000010000000000000000,
    22'b0000001001011100001010,
    22'b0000000010111000010100,
    22'b1111111111110101110001,
    22'b1111111100111101011100,
    22'b1111111010001111010111,
    22'b1111110111100001010010,
    22'b1111110011101011100001,
    22'b1111110001011100001010,
    22'b1111101111010111000011,
    22'b1111101100110011001101,
    22'b1111101000010100011111,
    22'b1111100100011110101110,
    22'b1111100000010100011111,
    22'b1111011100110011001101,
    22'b1111011010001111010111,
    22'b1111011000011110101110,
    22'b1111011000110011001101,
    22'b1111011001111010111000,
    22'b1111011100000000000000,
    22'b1111011100111101011100,
    22'b1111011011010111000011,
    22'b1111011011000010100100,
    22'b1111011011100001010010,
    22'b1111011101000111101100,
    22'b1111011110100011110110,
    22'b1111011110101110000101,
    22'b1111100001011100001010,
    22'b1111100100010100011111,
    22'b1111100110001111010111,
    22'b1111101000011110101110,
    22'b1111101110001111010111,
    22'b1111110000011110101110,
    22'b1111110010011001100110,
    22'b1111111000011110101110,
    22'b1111111111110101110001,
    22'b0000000100111101011100,
    22'b0000000011001100110011,
    22'b0000000011000010100100,
    22'b0000000000111101011100,
    22'b0000001101011100001010,
    22'b0000001001110000101001,
    22'b0000000011001100110011,
    22'b1111111011001100110011,
    22'b1111110101011100001010,
    22'b1111110101010001111011,
    22'b1111110100111101011100,
    22'b1111110010011001100110,
    22'b1111101011101011100001,
    22'b1111101010000101001000,
    22'b1111101011010111000011,
    22'b1111101100011110101110,
    22'b1111101101100110011010,
    22'b1111101110001111010111,
    22'b1111101101110000101001,
    22'b1111101100010100011111,
    22'b1111101010101110000101,
    22'b1111101001000111101100,
    22'b1111100111101011100001,
    22'b1111100110100011110110,
    22'b1111100110000101001000,
    22'b1111100110011001100110,
    22'b1111100111000010100100,
    22'b1111101000101000111101,
    22'b1111101001111010111000,
    22'b1111101011001100110011,
    22'b1111101100011110101110,
    22'b1111101101011100001010,
    22'b1111101111000010100100,
    22'b1111110001110000101001,
    22'b1111110101011100001010,
    22'b1111111000101000111101,
    22'b1111111111100001010010,
    22'b0000000100110011001101,
    22'b0000001100001010001111,
    22'b0000010101110000101001,
    22'b0000011100111101011100,
    22'b0000100001010001111011,
    22'b0000100100001010001111,
    22'b0000101011001100110011,
    22'b0000101111110101110001,
    22'b0000110000010100011111,
    22'b0000110001010001111011,
    22'b0000101111000010100100,
    22'b0000101110001111010111,
    22'b0000101101000111101100,
    22'b0000101000111101011100,
    22'b0000101000001010001111,
    22'b0000100111101011100001,
    22'b0000101000011110101110,
    22'b0000101011000010100100,
    22'b0000101111001100110011,
    22'b0000110110101110000101,
    22'b0000111100110011001101,
    22'b0001000010101110000101,
    22'b0001000110011001100110,
    22'b0001001011000010100100,
    22'b0001001110111000010100,
    22'b0001010000111101011100,
    22'b0001010000101000111101,
    22'b0001001110100011110110,
    22'b0001001100001010001111,
    22'b0001001001111010111000,
    22'b0001001001100110011010,
    22'b0001001011000010100100,
    22'b0001001110000101001000,
    22'b0001010010100011110110,
    22'b0001010110000101001000,
    22'b0001010101110000101001,
    22'b0001010000001010001111,
    22'b0001001011001100110011,
    22'b0001000100000000000000,
    22'b0001000000110011001101,
    22'b0000111111100001010010,
    22'b0000111111100001010010,
    22'b0001000000010100011111,
    22'b0000111110101110000101,
    22'b0000111101000111101100,
    22'b0000111100010100011111,
    22'b0000111011001100110011,
    22'b0000111000110011001101,
    22'b0000110101110000101001,
    22'b0000110010100011110110,
    22'b0000110000000000000000,
    22'b0000101101000111101100,
    22'b0000101011100001010010,
    22'b0000101100001010001111,
    22'b0000101110111000010100,
    22'b0000110010101110000101,
    22'b0000111010011001100110,
    22'b0001000000111101011100,
    22'b0001000110011001100110,
    22'b0001001010111000010100,
    22'b0001001101010001111011,
    22'b0001001110100011110110,
    22'b0001001011101011100001,
    22'b0001000111000010100100,
    22'b0001000001111010111000,
    22'b0000111010101110000101,
    22'b0000110101011100001010,
    22'b0000101111010111000011,
    22'b0000101000011110101110,
    22'b0000100010000101001000,
    22'b0000011010000101001000,
    22'b0000010100101000111101,
    22'b0000010000101000111101,
    22'b0000001101100110011010,
    22'b0000001011000010100100,
    22'b0000001010001111010111,
    22'b0000001010111000010100,
    22'b0000001100101000111101,
    22'b0000010000101000111101,
    22'b0000010100110011001101,
    22'b0000011001010001111011,
    22'b0000011101110000101001,
    22'b0000100001111010111000,
    22'b0000100110001111010111,
    22'b0000101000001010001111,
    22'b0000101000111101011100,
    22'b0000101000110011001101,
    22'b0000101000000000000000,
    22'b0000100111001100110011,
    22'b0000100110100011110110,
    22'b0000100101010001111011,
    22'b0000100011001100110011,
    22'b0000011111110101110001,
    22'b0000011100010100011111,
    22'b0000011011110101110001,
    22'b0000010100010100011111,
    22'b0000001001010001111011,
    22'b0000000011100001010010,
    22'b1111111101110000101001,
    22'b1111110111101011100001,
    22'b1111110001111010111000,
    22'b1111100101110000101001,
    22'b1111011110000101001000,
    22'b1111010110000101001000,
    22'b1111001000010100011111,
    22'b1110111001011100001010,
    22'b1110100000111101011100,
    22'b1101111010111000010100,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1110010101000111101100,
    22'b1110110111110101110001,
    22'b1111001100000000000000,
    22'b1111011011110101110001,
    22'b1111101010111000010100,
    22'b1111110101000111101100,
    22'b0000000100110011001101,
    22'b0000001101011100001010,
    22'b0000010010101110000101,
    22'b0000010101010001111011,
    22'b0000010101110000101001,
    22'b0000010011010111000011,
    22'b0000001110011001100110,
    22'b0000000111100001010010,
    22'b0000000000000000000000,
    22'b1111110110000101001000,
    22'b1111101111110101110001,
    22'b1111101010111000010100,
    22'b1111100111001100110011,
    22'b1111100100010100011111,
    22'b1111100000111101011100,
    22'b1111011111010111000011,
    22'b1111011101111010111000,
    22'b1111011100111101011100,
    22'b1111011100111101011100,
    22'b1111011101111010111000,
    22'b1111011110111000010100,
    22'b1111011111101011100001,
    22'b1111100000001010001111,
    22'b1111100001000111101100,
    22'b1111100010100011110110,
    22'b1111100011110101110001,
    22'b1111100110001111010111,
    22'b1111101000010100011111,
    22'b1111101010111000010100,
    22'b1111101100011110101110,
    22'b1111101110101110000101,
    22'b1111110000101000111101,
    22'b1111110011001100110011,
    22'b1111110101011100001010,
    22'b1111111000110011001101,
    22'b1111111111100001010010,
    22'b0000000101011100001010,
    22'b0000001011101011100001,
    22'b0000010010000101001000,
    22'b0000011001111010111000,
    22'b0000011111110101110001,
    22'b0000100101000111101100,
    22'b0000101001110000101001,
    22'b0000101111100001010010,
    22'b0000110011100001010010,
    22'b0000110111001100110011,
    22'b0000111010001111010111,
    22'b0000111100011110101110,
    22'b0000111101111010111000,
    22'b0000111110000101001000,
    22'b0000111101100110011010,
    22'b0000111100101000111101,
    22'b0000111011001100110011,
    22'b0000111010001111010111,
    22'b0000111001011100001010,
    22'b0000111000111101011100,
    22'b0000111000110011001101,
    22'b0000111000111101011100,
    22'b0000111000110011001101,
    22'b0000111000010100011111,
    22'b0000110111100001010010,
    22'b0000110110101110000101,
    22'b0000110110100011110110,
    22'b0000110111000010100100,
    22'b0000111000001010001111,
    22'b0000111001110000101001,
    22'b0000111011101011100001,
    22'b0000111100110011001101,
    22'b0000111101010001111011,
    22'b0000111101011100001010,
    22'b0000111100101000111101,
    22'b0000111011110101110001,
    22'b0000111011001100110011,
    22'b0000111010101110000101,
    22'b0000111010100011110110,
    22'b0000111010100011110110,
    22'b0000111010111000010100,
    22'b0000111011000010100100,
    22'b0000111010111000010100,
    22'b0000111010011001100110,
    22'b0000111010011001100110,
    22'b0000111010001111010111,
    22'b0000111000111101011100,
    22'b0000110110111000010100,
    22'b0000110101100110011010,
    22'b0000110100111101011100,
    22'b0000110101010001111011,
    22'b0000110100111101011100,
    22'b0000110011000010100100,
    22'b0000110001110000101001,
    22'b0000110000110011001101,
    22'b0000110000110011001101,
    22'b0000101110001111010111,
    22'b0000101100111101011100,
    22'b0000101100001010001111,
    22'b0000101100010100011111,
    22'b0000110100001010001111,
    22'b0000110101011100001010,
    22'b0000110001111010111000,
    22'b0000101101011100001010,
    22'b0000101011110101110001,
    22'b0000101001100110011010,
    22'b0000100110100011110110,
    22'b0000100010111000010100,
    22'b0000011101111010111000,
    22'b0000011011010111000011,
    22'b0000011001010001111011,
    22'b0000011000000000000000,
    22'b0000010111100001010010,
    22'b0000010111101011100001,
    22'b0000011000011110101110,
    22'b0000011001011100001010,
    22'b0000011010100011110110,
    22'b0000011100010100011111,
    22'b0000011101011100001010,
    22'b0000011110000101001000,
    22'b0000011110100011110110,
    22'b0000011110100011110110,
    22'b0000011110001111010111,
    22'b0000011101110000101001,
    22'b0000011101000111101100,
    22'b0000011100101000111101,
    22'b0000011100011110101110,
    22'b0000011100101000111101,
    22'b0000011100101000111101,
    22'b0000011100101000111101,
    22'b0000011100000000000000,
    22'b0000011011000010100100,
    22'b0000011001100110011010,
    22'b0000010111010111000011,
    22'b0000010101010001111011,
    22'b0000010010111000010100,
    22'b0000010000001010001111,
    22'b0000001100001010001111,
    22'b0000001001010001111011,
    22'b0000000110000101001000,
    22'b0000000010111000010100,
    22'b1111111110111000010100,
    22'b1111111011101011100001,
    22'b1111111000010100011111,
    22'b1111110100111101011100,
    22'b1111110000000000000000,
    22'b1111101100000000000000,
    22'b1111100111100001010010,
    22'b1111100001111010111000,
    22'b1111011000110011001101,
    22'b1111010000101000111101,
    22'b1111000111101011100001,
    22'b1110111110111000010100,
    22'b1110110011110101110001,
    22'b1110101100010100011111,
    22'b1110101001110000101001,
    22'b1110101011001100110011,
    22'b1110100110001111010111,
    22'b1110100000101000111101,
    22'b1110011011000010100100,
    22'b1110010101000111101100,
    22'b1110001101010001111011,
    22'b1110000111010111000011,
    22'b1110000000111101011100,
    22'b1101111010100011110110,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101111001000111101100,
    22'b1110000001000111101100,
    22'b1110001001010001111011,
    22'b1110010100010100011111,
    22'b1110011100011110101110,
    22'b1110100100000000000000,
    22'b1110101010011001100110,
    22'b1110110001010001111011,
    22'b1110110100111101011100,
    22'b1110110111001100110011,
    22'b1110110111110101110001,
    22'b1110110111000010100100,
    22'b1110110101100110011010,
    22'b1110110100000000000000,
    22'b1110110010000101001000,
    22'b1110110001010001111011,
    22'b1110110000111101011100,
    22'b1110110001000111101100,
    22'b1110110010001111010111,
    22'b1110110011100001010010,
    22'b1110110101000111101100,
    22'b1110110110011001100110,
    22'b1110111000010100011111,
    22'b1110111101000111101100,
    22'b1110111110101110000101,
    22'b1110111110001111010111,
    22'b1110111001111010111000,
    22'b1110110001000111101100,
    22'b1110100101010001111011,
    22'b1110011000001010001111,
    22'b1110001001000111101100,
    22'b1101111111110101110001,
    22'b1101110101100110011010,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100011110101110,
    22'b1101111000011110101110,
    22'b1101111100110011001101,
    22'b1110000100000000000000,
    22'b1110001001111010111000,
    22'b1110010000101000111101,
    22'b1110010110001111010111,
    22'b1110011101110000101001,
    22'b1110101111101011100001,
    22'b1110110010111000010100,
    22'b1110110101011100001010,
    22'b1110110101011100001010,
    22'b1110110011101011100001,
    22'b1110110000111101011100,
    22'b1110101011100001010010,
    22'b1110100111000010100100,
    22'b1110100010101110000101,
    22'b1110011110001111010111,
    22'b1110011100001010001111,
    22'b1110011011110101110001,
    22'b1110011101010001111011,
    22'b1110100001010001111011,
    22'b1110100101011100001010,
    22'b1110101010001111010111,
    22'b1110101111010111000011,
    22'b1110110110000101001000,
    22'b1110111010100011110110,
    22'b1110111101110000101001,
    22'b1111000000101000111101,
    22'b1111000001011100001010,
    22'b1111000000001010001111,
    22'b1110111100011110101110,
    22'b1110110101000111101100,
    22'b1110110000001010001111,
    22'b1110101101000111101100,
    22'b1110101011110101110001,
    22'b1110101100011110101110,
    22'b1110101110011001100110,
    22'b1110110000111101011100,
    22'b1110110101011100001010,
    22'b1110111000111101011100,
    22'b1110111100010100011111,
    22'b1110111111001100110011,
    22'b1111000010111000010100,
    22'b1111000101100110011010,
    22'b1111001000110011001101,
    22'b1111001110000101001000,
    22'b1111010010101110000101,
    22'b1111100110111000010100,
    22'b1111101010101110000101,
    22'b1111101101000111101100,
    22'b1111101110111000010100,
    22'b1111110000011110101110,
    22'b1111110010011001100110,
    22'b1111110011110101110001,
    22'b1111110100111101011100,
    22'b1111110100110011001101,
    22'b1111110100001010001111,
    22'b1111110011010111000011,
    22'b1111110010011001100110,
    22'b1111110001011100001010,
    22'b1111110001000111101100,
    22'b1111110001000111101100,
    22'b1111110001010001111011,
    22'b1111110001010001111011,
    22'b1111110001010001111011,
    22'b1111110000111101011100,
    22'b1111110000101000111101,
    22'b1111110000011110101110,
    22'b1111110000110011001101,
    22'b1111110001100110011010,
    22'b1111110011000010100100,
    22'b1111110100001010001111,
    22'b1111110101010001111011,
    22'b1111110110100011110110,
    22'b1111111000110011001101,
    22'b1111111010111000010100,
    22'b1111111101011100001010,
    22'b0000000000101000111101,
    22'b0000000101100110011010,
    22'b0000011011001100110011,
    22'b0000100001000111101100,
    22'b0000101010000101001000,
    22'b0000110001110000101001,
    22'b0000111010011001100110,
    22'b0001000111101011100001,
    22'b0001010010100011110110,
    22'b0001011101110000101001,
    22'b0001011001100110011010,
    22'b0001001100011110101110,
    22'b0001001000001010001111,
    22'b0001001000011110101110,
    22'b0001001100011110101110,
    22'b0001010100010100011111,
    22'b0001011100010100011111,
    22'b0001100100110011001101,
    22'b0001110011000010100100,
    22'b0001111110100011110110,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0001111001100110011010,
    22'b0001101011001100110011,
    22'b0001100001010001111011,
    22'b0001011010111000010100,
    22'b0001011010100011110110,
    22'b0001011101010001111011,
    22'b0001100010001111010111,
    22'b0001101010111000010100,
    22'b0001110010000101001000,
    22'b0001111001000111101100,
    22'b0001111111000010100100,
    22'b0010000101010001111011,
    22'b0010001000000000000000,
    22'b0010001000110011001101,
    22'b0010000111001100110011,
    22'b0010000101000111101100,
    22'b0010000010111000010100,
    22'b0010000001100110011010,
    22'b0010000001100110011010,
    22'b0010000010011001100110,
    22'b0010000100001010001111,
    22'b0010000110111000010100,
    22'b0010001010101110000101,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011001100110011,
    22'b0010001010000101001000,
    22'b0010001001010001111011,
    22'b0010001001100110011010,
    22'b0010001010011001100110,
    22'b0010001011001100110011,
    22'b0010001010100011110110,
    22'b0010001000001010001111,
    22'b0010000101000111101100,
    22'b0010000001100110011010,
    22'b0001111101111010111000,
    22'b0001111010011001100110,
    22'b0001110110011001100110,
    22'b0001110100000000000000,
    22'b0001110010000101001000,
    22'b0001110000110011001101,
    22'b0001101111100001010010,
    22'b0001101110100011110110,
    22'b0001101101100110011010,
    22'b0001101100110011001101,
    22'b0001101011001100110011,
    22'b0001101001111010111000,
    22'b0001101000000000000000,
    22'b0001100101111010111000,
    22'b0001100010111000010100,
    22'b0001100000110011001101,
    22'b0001011110111000010100,
    22'b0001011101110000101001,
    22'b0001011100001010001111,
    22'b0001011010001111010111,
    22'b0001010111101011100001,
    22'b0001010100101000111101,
    22'b0001010001010001111011,
    22'b0001001110111000010100,
    22'b0001001110011001100110,
    22'b0001001110011001100110,
    22'b0001001001011100001010,
    22'b0001000100001010001111,
    22'b0001000000110011001101,
    22'b0001000010100011110110,
    22'b0001001001000111101100,
    22'b0001001101011100001010,
    22'b0001001111001100110011,
    22'b0001010000001010001111,
    22'b0001010000110011001101,
    22'b0001010001000111101100,
    22'b0001010000010100011111,
    22'b0001010000011110101110,
    22'b0001010001110000101001,
    22'b0001010010011001100110,
    22'b0001010010101110000101,
    22'b0001010010111000010100,
    22'b0001010011010111000011,
    22'b0001010100000000000000,
    22'b0001010100010100011111,
    22'b0001010011110101110001,
    22'b0001010010101110000101,
    22'b0001010000110011001101,
    22'b0001001111010111000011,
    22'b0001001101111010111000,
    22'b0001001100000000000000,
    22'b0001001001100110011010,
    22'b0001001000001010001111,
    22'b0001000110111000010100,
    22'b0001000100111101011100,
    22'b0001000001110000101001,
    22'b0000111110101110000101,
    22'b0000111011101011100001,
    22'b0000111010000101001000,
    22'b0000111010100011110110,
    22'b0000111010111000010100,
    22'b0000111001111010111000,
    22'b0000110110011001100110,
    22'b0000110100111101011100,
    22'b0000110010011001100110,
    22'b0000101111100001010010,
    22'b0000101100011110101110,
    22'b0000101010000101001000,
    22'b0000100111100001010010,
    22'b0000100101010001111011,
    22'b0000100011000010100100,
    22'b0000100001100110011010,
    22'b0000100000000000000000,
    22'b0000011110001111010111,
    22'b0000011100010100011111,
    22'b0000011011001100110011,
    22'b0000011001100110011010,
    22'b0000010111110101110001,
    22'b0000010100101000111101,
    22'b0000010001100110011010,
    22'b0000001101110000101001,
    22'b0000001010001111010111,
    22'b0000000110011001100110,
    22'b0000000011101011100001,
    22'b0000000001000111101100,
    22'b1111111110101110000101,
    22'b1111111011110101110001,
    22'b1111111001111010111000,
    22'b1111111000011110101110,
    22'b1111110111010111000011,
    22'b1111110110011001100110,
    22'b1111110101110000101001,
    22'b1111110100111101011100,
    22'b1111110011010111000011,
    22'b1111110001110000101001,
    22'b1111110000001010001111,
    22'b1111101110111000010100,
    22'b1111101101011100001010,
    22'b1111101101100110011010,
    22'b1111101101010001111011,
    22'b1111101101011100001010,
    22'b1111101101110000101001,
    22'b1111101110111000010100,
    22'b1111110000001010001111,
    22'b1111110010101110000101,
    22'b1111110011100001010010,
    22'b1111110101010001111011,
    22'b1111110101100110011010,
    22'b1111110110101110000101,
    22'b1111110110000101001000,
    22'b1111110101100110011010,
    22'b1111110101000111101100,
    22'b1111110110100011110110,
    22'b1111110110011001100110,
    22'b1111110110001111010111,
    22'b1111110101011100001010,
    22'b1111110100001010001111,
    22'b1111110010101110000101,
    22'b1111110001011100001010,
    22'b1111110000010100011111,
    22'b1111101111010111000011,
    22'b1111101110001111010111,
    22'b1111101100110011001101,
    22'b1111101010100011110110,
    22'b1111101000101000111101,
    22'b1111100111000010100100,
    22'b1111011110111000010100,
    22'b1111011100101000111101,
    22'b1111011001100110011010,
    22'b1111010110000101001000,
    22'b1111010000010100011111,
    22'b1111001011101011100001,
    22'b1111000110100011110110,
    22'b1110111111001100110011,
    22'b1110111001100110011010,
    22'b1110110100101000111101,
    22'b1110110000011110101110,
    22'b1110101010000101001000,
    22'b1110100110100011110110,
    22'b1110100011101011100001,
    22'b1110100010111000010100,
    22'b1110100011110101110001,
    22'b1110100110001111010111,
    22'b1110101010001111010111,
    22'b1110101110101110000101,
    22'b1110110101010001111011,
    22'b1110111001111010111000,
    22'b1110111101011100001010,
    22'b1110111111110101110001,
    22'b1111000001111010111000,
    22'b1111000010100011110110,
    22'b1111000010001111010111,
    22'b1111000000011110101110,
    22'b1110111011001100110011,
    22'b1110110110000101001000,
    22'b1110110000101000111101,
    22'b1110101010101110000101,
    22'b1110100111100001010010,
    22'b1110100101010001111011,
    22'b1110100100000000000000,
    22'b1110100011001100110011,
    22'b1110100011001100110011,
    22'b1110100011000010100100,
    22'b1110100011000010100100,
    22'b1110100011010111000011,
    22'b1110100100001010001111,
    22'b1110100101000111101100,
    22'b1110100110000101001000,
    22'b1110100111010111000011,
    22'b1110100111110101110001,
    22'b1110100111110101110001,
    22'b1110100111101011100001,
    22'b1110100111100001010010,
    22'b1110100111001100110011,
    22'b1110100110000101001000,
    22'b1110100100011110101110,
    22'b1110100001100110011010,
    22'b1110011111001100110011,
    22'b1110011100110011001101,
    22'b1110011010100011110110,
    22'b1110011000110011001101,
    22'b1110010111001100110011,
    22'b1110010110111000010100,
    22'b1110010111001100110011,
    22'b1110011000000000000000,
    22'b1110011001011100001010,
    22'b1110011010000101001000,
    22'b1110011010101110000101,
    22'b1110011011001100110011,
    22'b1110011011100001010010,
    22'b1110011100101000111101,
    22'b1110011110011001100110,
    22'b1110100000111101011100,
    22'b1110100100001010001111,
    22'b1110101000011110101110,
    22'b1110101010111000010100,
    22'b1110101100011110101110,
    22'b1110101100101000111101,
    22'b1110101011101011100001,
    22'b1110001011110101110001,
    22'b1110000101000111101100,
    22'b1101111111001100110011,
    22'b1101111001010001111011,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101111010111000010100,
    22'b1110000001111010111000,
    22'b1110001000110011001101,
    22'b1110010001011100001010,
    22'b1110010111001100110011,
    22'b1110011100011110101110,
    22'b1110100000111101011100,
    22'b1110100101011100001010,
    22'b1110100111010111000011,
    22'b1110101000101000111101,
    22'b1110101000110011001101,
    22'b1110100111101011100001,
    22'b1110100101011100001010,
    22'b1110100010001111010111,
    22'b1110011101110000101001,
    22'b1110010110000101001000,
    22'b1110001111100001010010,
    22'b1110001000110011001101,
    22'b1110000010100011110110,
    22'b1101111100000000000000,
    22'b1101111000101000111101,
    22'b1101110110111000010100,
    22'b1101110110111000010100,
    22'b1101111000110011001101,
    22'b1101111011101011100001,
    22'b1101111111000010100100,
    22'b1110000010111000010100,
    22'b1110000111101011100001,
    22'b1110001010101110000101,
    22'b1110001100101000111101,
    22'b1110001101010001111011,
    22'b1110001100001010001111,
    22'b1110001010100011110110,
    22'b1110001000011110101110,
    22'b1110000110001111010111,
    22'b1110000011010111000011,
    22'b1110000001110000101001,
    22'b1110000001010001111011,
    22'b1110000100111101011100,
    22'b1110000111100001010010,
    22'b1110001010011001100110,
    22'b1110001101000111101100,
    22'b1110010001010001111011,
    22'b1110010100101000111101,
    22'b1110011000010100011111,
    22'b1110011100000000000000,
    22'b1110100000010100011111,
    22'b1110100010011001100110,
    22'b1110100011110101110001,
    22'b1110100100001010001111,
    22'b1110100011110101110001,
    22'b1110100010011001100110,
    22'b1110100001010001111011,
    22'b1110011111000010100100,
    22'b1110011100010100011111,
    22'b1110011000010100011111,
    22'b1110010101000111101100,
    22'b1110010010011001100110,
    22'b1110010000000000000000,
    22'b1110001101110000101001,
    22'b1110001100101000111101,
    22'b1110001100001010001111,
    22'b1110001100010100011111,
    22'b1110001100110011001101,
    22'b1110001101100110011010,
    22'b1110001110100011110110,
    22'b1110001111110101110001,
    22'b1110010000111101011100,
    22'b1110010010000101001000,
    22'b1110010011101011100001,
    22'b1110010110001111010111,
    22'b1110011000111101011100,
    22'b1110011011101011100001,
    22'b1110011110101110000101,
    22'b1110100010100011110110,
    22'b1110100101010001111011,
    22'b1110100111110101110001,
    22'b1110101010001111010111,
    22'b1110101101000111101100,
    22'b1110101111001100110011,
    22'b1110110001010001111011,
    22'b1110110011100001010010,
    22'b1110110110101110000101,
    22'b1110111001011100001010,
    22'b1110111100001010001111,
    22'b1110111111000010100100,
    22'b1111001000111101011100,
    22'b1111001000111101011100,
    22'b1111000111010111000011,
    22'b1111000111001100110011,
    22'b1111001010100011110110,
    22'b1111001100110011001101,
    22'b1111010001110000101001,
    22'b1111100000101000111101,
    22'b1111101101000111101100,
    22'b0000001100000000000000,
    22'b0000110000111101011100,
    22'b0000110010100011110110,
    22'b0000001100010100011111,
    22'b1111110100001010001111,
    22'b1111011111100001010010,
    22'b1111010010111000010100,
    22'b1111001110111000010100,
    22'b1111001111010111000011,
    22'b1111010010100011110110,
    22'b1111010111100001010010,
    22'b1111011011101011100001,
    22'b1111100000000000000000,
    22'b1111100101000111101100,
    22'b1111101000011110101110,
    22'b1111101011010111000011,
    22'b1111101101111010111000,
    22'b1111110001011100001010,
    22'b1111110100010100011111,
    22'b1111110111010111000011,
    22'b1111111010011001100110,
    22'b1111111110001111010111,
    22'b0000000000111101011100,
    22'b0000000011010111000011,
    22'b0000000101110000101001,
    22'b0000001000010100011111,
    22'b0000001001111010111000,
    22'b0000001011010111000011,
    22'b0000001100111101011100,
    22'b0000010110100011110110,
    22'b0000011000011110101110,
    22'b0000011010000101001000,
    22'b0000011011100001010010,
    22'b0000011100000000000000,
    22'b0000011100010100011111,
    22'b0000011100000000000000,
    22'b0000011011000010100100,
    22'b0000011010001111010111,
    22'b0000011001011100001010,
    22'b0000011000011110101110,
    22'b0000010111000010100100,
    22'b0000010101100110011010,
    22'b0000010100001010001111,
    22'b0000010010111000010100,
    22'b0000010001010001111011,
    22'b0000010000101000111101,
    22'b0000010000101000111101,
    22'b0000010000110011001101,
    22'b0000010001100110011010,
    22'b0000010010111000010100,
    22'b0000010100101000111101,
    22'b0000010111000010100100,
    22'b0000011011010111000011,
    22'b0000011111000010100100,
    22'b0000100011001100110011,
    22'b0000101000000000000000,
    22'b0000101111001100110011,
    22'b0000110100101000111101,
    22'b0000111010011001100110,
    22'b0001000011000010100100,
    22'b0001001001100110011010,
    22'b0001010000101000111101,
    22'b0001010111110101110001,
    22'b0001100001111010111000,
    22'b0001101001100110011010,
    22'b0001110001011100001010,
    22'b0001111001011100001010,
    22'b0010000100001010001111,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010000101011100001010,
    22'b0001111011000010100100,
    22'b0001110001000111101100,
    22'b0001101000011110101110,
    22'b0001100000111101011100,
    22'b0001011001011100001010,
    22'b0001010101110000101001,
    22'b0001010011101011100001,
    22'b0001010010111000010100,
    22'b0001010010101110000101,
    22'b0001010011100001010010,
    22'b0001010100011110101110,
    22'b0001010101000111101100,
    22'b0001010101110000101001,
    22'b0001010110001111010111,
    22'b0001010110000101001000,
    22'b0001010101110000101001,
    22'b0001010110011001100110,
    22'b0001010111100001010010,
    22'b0001011001010001111011,
    22'b0001011010001111010111,
    22'b0001011011100001010010,
    22'b0001011100110011001101,
    22'b0001011101110000101001,
    22'b0001011111110101110001,
    22'b0001100000111101011100,
    22'b0001100001100110011010,
    22'b0001100010111000010100,
    22'b0001100100111101011100,
    22'b0001100110011001100110,
    22'b0001100111100001010010,
    22'b0001101000110011001101,
    22'b0001101001111010111000,
    22'b0001101001111010111000,
    22'b0001101001011100001010,
    22'b0001101000011110101110,
    22'b0001100110111000010100,
    22'b0001100100101000111101,
    22'b0001100010000101001000,
    22'b0001011111001100110011,
    22'b0001011100000000000000,
    22'b0001011000000000000000,
    22'b0001010000110011001101,
    22'b0001001011110101110001,
    22'b0001000110111000010100,
    22'b0001000010000101001000,
    22'b0000111100011110101110,
    22'b0000111000011110101110,
    22'b0000110100101000111101,
    22'b0000110001110000101001,
    22'b0000101111101011100001,
    22'b0000101110000101001000,
    22'b0000101101010001111011,
    22'b0000101101010001111011,
    22'b0000101101100110011010,
    22'b0000101110101110000101,
    22'b0000110000001010001111,
    22'b0000110001111010111000,
    22'b0000110011010111000011,
    22'b0000110100010100011111,
    22'b0000110100110011001101,
    22'b0000110101000111101100,
    22'b0000110101011100001010,
    22'b0000110111000010100100,
    22'b0000110110101110000101,
    22'b0000110011001100110011,
    22'b0000110000101000111101,
    22'b0000101110111000010100,
    22'b0000101101100110011010,
    22'b0000101100000000000000,
    22'b0000101010011001100110,
    22'b0000101000011110101110,
    22'b0000100110101110000101,
    22'b0000100101000111101100,
    22'b0000100010111000010100,
    22'b0000100001000111101100,
    22'b0000011111101011100001,
    22'b0000011110101110000101,
    22'b0000011110011001100110,
    22'b0000011110111000010100,
    22'b0000011110000101001000,
    22'b0000011000111101011100,
    22'b0000001100110011001101,
    22'b0000000111100001010010,
    22'b0000000000010100011111,
    22'b1111111000011110101110,
    22'b1111110000010100011111,
    22'b1111101101000111101100,
    22'b1111101110001111010111,
    22'b1111110011100001010010,
    22'b1111111010011001100110,
    22'b0000000001110000101001,
    22'b0000001000000000000000,
    22'b0000001111000010100100,
    22'b0000010101110000101001,
    22'b0000011100111101011100,
    22'b0000100110100011110110,
    22'b0000101101100110011010,
    22'b0000110100001010001111,
    22'b0000111001110000101001,
    22'b0000111111001100110011,
    22'b0001000001110000101001,
    22'b0001000011010111000011,
    22'b0001000100000000000000,
    22'b0001000100001010001111,
    22'b0001000011110101110001,
    22'b0001000011010111000011,
    22'b0001000010111000010100,
    22'b0001000010000101001000,
    22'b0001000000101000111101,
    22'b0000111101100110011010,
    22'b0000111000111101011100,
    22'b0000110010101110000101,
    22'b0000101100001010001111,
    22'b0000100100000000000000,
    22'b0000011111101011100001,
    22'b0000011100101000111101,
    22'b0000011010100011110110,
    22'b0000011001010001111011,
    22'b0000010111100001010010,
    22'b0000010101111010111000,
    22'b0000010011101011100001,
    22'b0000010001000111101100,
    22'b0000001101010001111011,
    22'b0000001010100011110110,
    22'b0000001000011110101110,
    22'b0000000110101110000101,
    22'b0000000101011100001010,
    22'b0000000100010100011111,
    22'b0000000011101011100001,
    22'b0000000011001100110011,
    22'b0000000010101110000101,
    22'b0000000010100011110110,
    22'b0000000010100011110110,
    22'b0000000011101011100001,
    22'b0000001101010001111011,
    22'b0000010100101000111101,
    22'b0000011011101011100001,
    22'b0000011101100110011010,
    22'b0000011111000010100100,
    22'b0000011111100001010010,
    22'b0000011110100011110110,
    22'b0000011100010100011111,
    22'b0000011001010001111011,
    22'b0000010101000111101100,
    22'b0000010010001111010111,
    22'b0000001111110101110001,
    22'b0000001101100110011010,
    22'b0000001011100001010010,
    22'b0000001000101000111101,
    22'b0000000110011001100110,
    22'b0000000011101011100001,
    22'b0000000000110011001101,
    22'b1111111100101000111101,
    22'b1111111001011100001010,
    22'b1111110110011001100110,
    22'b1111110011010111000011,
    22'b1111101111010111000011,
    22'b1111101100010100011111,
    22'b1111101001011100001010,
    22'b1111100110101110000101,
    22'b1111100100000000000000,
    22'b1111100000001010001111,
    22'b1111011101000111101100,
    22'b1111011001111010111000,
    22'b1111010110001111010111,
    22'b1111010001110000101001,
    22'b1111001110101110000101,
    22'b1111001100001010001111,
    22'b1111001010100011110110,
    22'b1111001001010001111011,
    22'b1111001001010001111011,
    22'b1111001001111010111000,
    22'b1111001010111000010100,
    22'b1111001100111101011100,
    22'b1111001110100011110110,
    22'b1111010000001010001111,
    22'b1111010001100110011010,
    22'b1111010011101011100001,
    22'b1111010101000111101100,
    22'b1111010110101110000101,
    22'b1111011000010100011111,
    22'b1111011010001111010111,
    22'b1111011011001100110011,
    22'b1111011100000000000000,
    22'b1111011100110011001101,
    22'b1111011101100110011010,
    22'b1111011111000010100100,
    22'b1111100000010100011111,
    22'b1111100001110000101001,
    22'b1111100011000010100100,
    22'b1111100100011110101110,
    22'b1111100101011100001010,
    22'b1111100110000101001000,
    22'b1111100110100011110110,
    22'b1111100110111000010100,
    22'b1111100110111000010100,
    22'b1111100110111000010100,
    22'b1111100110101110000101,
    22'b1111100110101110000101,
    22'b1111100110101110000101,
    22'b1111100111000010100100,
    22'b1111100111001100110011,
    22'b1111100111100001010010,
    22'b1111101000000000000000,
    22'b1111101000001010001111,
    22'b1111100111110101110001,
    22'b1111100111100001010010,
    22'b1111100110111000010100,
    22'b1111100110011001100110,
    22'b1111100101111010111000,
    22'b1111100101110000101001,
    22'b1111100101110000101001,
    22'b1111100101111010111000,
    22'b1111100101111010111000,
    22'b1111100110100011110110,
    22'b1111100111000010100100,
    22'b1111100111100001010010,
    22'b1111100111110101110001,
    22'b1111100111110101110001,
    22'b1111100111100001010010,
    22'b1111100111001100110011,
    22'b1111100110111000010100,
    22'b1111100110100011110110,
    22'b1111100110100011110110,
    22'b1111100110100011110110,
    22'b1111100110101110000101,
    22'b1111100111001100110011,
    22'b1111101000000000000000,
    22'b1111101001010001111011,
    22'b1111101010101110000101,
    22'b1111101100111101011100,
    22'b1111101110011001100110,
    22'b1111101111100001010010,
    22'b1111110000101000111101,
    22'b1111110001111010111000,
    22'b1111110010111000010100,
    22'b1111110011110101110001,
    22'b1111110100110011001101,
    22'b1111110101011100001010,
    22'b1111110101110000101001,
    22'b1111110110000101001000,
    22'b1111110110000101001000,
    22'b1111110101111010111000,
    22'b1111110101110000101001,
    22'b1111110101011100001010,
    22'b1111110100111101011100,
    22'b1111110100011110101110,
    22'b1111110011101011100001,
    22'b1111110010111000010100,
    22'b1111110001111010111000,
    22'b1111110000111101011100,
    22'b1111110000000000000000,
    22'b1111101110000101001000,
    22'b1111101010111000010100,
    22'b1111101001010001111011,
    22'b1111101000110011001101,
    22'b1111101000110011001101,
    22'b1111101000110011001101,
    22'b1111101000111101011100,
    22'b1111101000110011001101,
    22'b1111101001000111101100,
    22'b1111101001111010111000,
    22'b1111101011000010100100,
    22'b1111101100010100011111,
    22'b1111101101010001111011,
    22'b1111101101011100001010,
    22'b1111101101100110011010,
    22'b1111101101110000101001,
    22'b1111101101100110011010,
    22'b1111101101011100001010,
    22'b1111101101010001111011,
    22'b1111101100110011001101,
    22'b1111101100011110101110,
    22'b1111101100010100011111,
    22'b1111101100001010001111,
    22'b1111101011110101110001,
    22'b1111101011110101110001,
    22'b1111101011110101110001,
    22'b1111101100000000000000,
    22'b1111101100010100011111,
    22'b1111101100011110101110,
    22'b1111101100101000111101,
    22'b1111101100111101011100,
    22'b1111101100111101011100,
    22'b1111101101000111101100,
    22'b1111101101000111101100,
    22'b1111101101010001111011,
    22'b1111101101010001111011,
    22'b1111101101000111101100,
    22'b1111101011001100110011,
    22'b1111101010111000010100,
    22'b1111101010100011110110,
    22'b1111101001111010111000,
    22'b1111101001010001111011,
    22'b1111101000011110101110,
    22'b1111100111100001010010,
    22'b1111100110101110000101,
    22'b1111100110000101001000,
    22'b1111100101000111101100,
    22'b1111100100001010001111,
    22'b1111100010011001100110,
    22'b1111100001010001111011,
    22'b1111100000010100011111,
    22'b1111011111100001010010,
    22'b1111011111001100110011,
    22'b1111011111000010100100,
    22'b1111011110111000010100,
    22'b1111011111000010100100,
    22'b1111011111001100110011,
    22'b1111011111101011100001,
    22'b1111100000101000111101,
    22'b1111100001110000101001,
    22'b1111100011000010100100,
    22'b1111100100010100011111,
    22'b1111100101111010111000,
    22'b1111100111000010100100,
    22'b1111101000001010001111,
    22'b1111101001000111101100,
    22'b1111101010000101001000,
    22'b1111101010001111010111,
    22'b1111101010011001100110,
    22'b1111101011000010100100,
    22'b1111101011101011100001,
    22'b1111101100011110101110,
    22'b1111101101100110011010,
    22'b1111101110001111010111,
    22'b1111101111000010100100,
    22'b1111101111101011100001,
    22'b1111110000101000111101,
    22'b1111110001010001111011,
    22'b1111110001111010111000,
    22'b1111110010100011110110,
    22'b1111110011010111000011,
    22'b1111110011101011100001,
    22'b1111110011110101110001,
    22'b1111110100000000000000,
    22'b1111110100000000000000,
    22'b1111110011110101110001,
    22'b1111110011110101110001,
    22'b1111110100000000000000,
    22'b1111110100001010001111,
    22'b1111110100010100011111,
    22'b1111110100110011001101,
    22'b1111110101010001111011,
    22'b1111110101110000101001,
    22'b1111110110011001100110,
    22'b1111110110111000010100,
    22'b1111110111000010100100,
    22'b1111110110111000010100,
    22'b1111110110011001100110,
    22'b1111110101100110011010,
    22'b1111110000011110101110,
    22'b1111101110001111010111,
    22'b1111101011101011100001,
    22'b1111101010011001100110,
    22'b1111101001100110011010,
    22'b1111101001000111101100,
    22'b1111101001010001111011,
    22'b1111101001110000101001,
    22'b1111101010000101001000,
    22'b1111101010100011110110,
    22'b1111101010111000010100,
    22'b1111101011001100110011,
    22'b1111101011101011100001,
    22'b1111101100011110101110,
    22'b1111101101011100001010,
    22'b1111101110100011110110,
    22'b1111110000010100011111,
    22'b1111110001110000101001,
    22'b1111110011001100110011,
    22'b1111110100110011001101,
    22'b1111110110101110000101,
    22'b1111111000000000000000,
    22'b1111111001010001111011,
    22'b1111111010100011110110,
    22'b1111111100011110101110,
    22'b1111111110001111010111,
    22'b0000000000001010001111,
    22'b0000000010101110000101,
    22'b0000000100010100011111,
    22'b0000000101100110011010,
    22'b0000000110101110000101,
    22'b0000001010100011110110,
    22'b0000001011010111000011,
    22'b0000001100000000000000,
    22'b0000001100111101011100,
    22'b0000001101110000101001,
    22'b0000001110100011110110,
    22'b0000001111010111000011,
    22'b0000001111110101110001,
    22'b0000010000000000000000,
    22'b0000001111110101110001,
    22'b0000001111100001010010,
    22'b0000001111001100110011,
    22'b0000001110111000010100,
    22'b0000001110100011110110,
    22'b0000001101111010111000,
    22'b0000001100111101011100,
    22'b0000001011110101110001,
    22'b0000001001100110011010,
    22'b0000000111100001010010,
    22'b0000000101010001111011,
    22'b0000000010101110000101,
    22'b1111111111101011100001,
    22'b1111111101100110011010,
    22'b1111111011101011100001,
    22'b1111111001111010111000,
    22'b1111111001000111101100,
    22'b1111111000101000111101,
    22'b1111111000101000111101,
    22'b1111111001000111101100,
    22'b1111111001100110011010,
    22'b1111111010001111010111,
    22'b1111111001011100001010,
    22'b1111111000010100011111,
    22'b1111110111000010100100,
    22'b1111110101100110011010,
    22'b1111110100110011001101,
    22'b1111110100010100011111,
    22'b1111110100000000000000,
    22'b1111110011100001010010,
    22'b1111110011000010100100,
    22'b1111110010111000010100,
    22'b1111110011000010100100,
    22'b1111110011101011100001,
    22'b1111110100000000000000,
    22'b1111110011110101110001,
    22'b1111110010111000010100,
    22'b1111110001100110011010,
    22'b1111110000011110101110,
    22'b1111101111100001010010,
    22'b1111101110101110000101,
    22'b1111101110101110000101,
    22'b1111101110101110000101,
    22'b1111101111010111000011,
    22'b1111110000000000000000,
    22'b1111110000110011001101,
    22'b1111110001111010111000,
    22'b1111110011001100110011,
    22'b1111110100010100011111,
    22'b1111110101011100001010,
    22'b1111110110011001100110,
    22'b1111110111001100110011,
    22'b1111110111001100110011,
    22'b1111110010111000010100,
    22'b1111110001000111101100,
    22'b1111101111110101110001,
    22'b1111101111000010100100,
    22'b1111101110001111010111,
    22'b1111101101111010111000,
    22'b1111101101110000101001,
    22'b1111101101111010111000,
    22'b1111101110001111010111,
    22'b1111101110001111010111,
    22'b1111101110011001100110,
    22'b1111101110001111010111,
    22'b1111101110000101001000,
    22'b1111101110000101001000,
    22'b1111101110011001100110,
    22'b1111101110101110000101,
    22'b1111101111010111000011,
    22'b1111101111101011100001,
    22'b1111101111101011100001,
    22'b1111101111010111000011,
    22'b1111101110111000010100,
    22'b1111101101111010111000,
    22'b1111101100101000111101,
    22'b1111101011000010100100,
    22'b1111101001111010111000,
    22'b1111101001000111101100,
    22'b1111101000001010001111,
    22'b1111100111100001010010,
    22'b1111100111110101110001,
    22'b1111101000010100011111,
    22'b1111101000000000000000,
    22'b1111100110101110000101,
    22'b1111100011100001010010,
    22'b1111100000101000111101,
    22'b1111011101110000101001,
    22'b1111011010101110000101,
    22'b1111010110101110000101,
    22'b1111010011001100110011,
    22'b1111001111110101110001,
    22'b1111001100101000111101,
    22'b1111001000110011001101,
    22'b1111000110111000010100,
    22'b1111000101111010111000,
    22'b1111000110011001100110,
    22'b1111001000001010001111,
    22'b1111001010100011110110,
    22'b1111001010011001100110,
    22'b1111001011010111000011,
    22'b1111001011110101110001,
    22'b1111001100010100011111,
    22'b1111001100000000000000,
    22'b1111001010101110000101,
    22'b1111001010001111010111,
    22'b1111001001111010111000,
    22'b1111001001011100001010,
    22'b1111001001110000101001,
    22'b1111001001111010111000,
    22'b1111001010101110000101,
    22'b1111010010001111010111,
    22'b1111010100001010001111,
    22'b1111010101110000101001,
    22'b1111010111000010100100,
    22'b1111010111010111000011,
    22'b1111011000001010001111,
    22'b1111011000111101011100,
    22'b1111011001111010111000,
    22'b1111011001010001111011,
    22'b1111011001000111101100,
    22'b1111011010000101001000,
    22'b1111011010101110000101,
    22'b1111011010101110000101,
    22'b1111011010000101001000,
    22'b1111011000011110101110,
    22'b1111010110011001100110,
    22'b1111010100110011001101,
    22'b1111010011100001010010,
    22'b1111010001100110011010,
    22'b1111001111001100110011,
    22'b1111001110100011110110,
    22'b1111001111001100110011,
    22'b1111010000110011001101,
    22'b1111010001110000101001,
    22'b1111010010001111010111,
    22'b1111010011000010100100,
    22'b1111010011100001010010,
    22'b1111010011110101110001,
    22'b1111010011010111000011,
    22'b1111010101000111101100,
    22'b1111011100110011001101,
    22'b1111011001100110011010,
    22'b1111010111100001010010,
    22'b1111010110101110000101,
    22'b1111010101100110011010,
    22'b1111010011000010100100,
    22'b1111010000111101011100,
    22'b1111010001010001111011,
    22'b1111010011110101110001,
    22'b1111010011001100110011,
    22'b1111010101000111101100,
    22'b1111010101110000101001,
    22'b1111010110001111010111,
    22'b1111010101110000101001,
    22'b1111010110000101001000,
    22'b1111011000010100011111,
    22'b1111010011101011100001,
    22'b1111010011001100110011,
    22'b1111010000000000000000,
    22'b1111010001011100001010,
    22'b1111010010001111010111,
    22'b1111010001000111101100,
    22'b1111010011101011100001,
    22'b1111010100111101011100,
    22'b1111011000111101011100,
    22'b1111011100011110101110,
    22'b1111100000010100011111,
    22'b1111100011100001010010,
    22'b1111100011100001010010,
    22'b1111100101110000101001,
    22'b1111101000011110101110,
    22'b1111110010000101001000,
    22'b1111110011010111000011,
    22'b1111110100011110101110,
    22'b1111110101100110011010,
    22'b1111110110011001100110,
    22'b1111110111001100110011,
    22'b1111111000000000000000,
    22'b1111111000111101011100,
    22'b1111111001110000101001,
    22'b1111111010101110000101,
    22'b1111111011101011100001,
    22'b1111111101010001111011,
    22'b1111111110001111010111,
    22'b1111111111001100110011,
    22'b1111111111110101110001,
    22'b0000000000101000111101,
    22'b0000000000111101011100,
    22'b0000000000101000111101,
    22'b1111111111100001010010,
    22'b1111111101110000101001,
    22'b1111111100101000111101,
    22'b1111111100000000000000,
    22'b1111111011101011100001,
    22'b1111111011101011100001,
    22'b1111111100000000000000,
    22'b1111111100011110101110,
    22'b1111111101000111101100,
    22'b1111111110000101001000,
    22'b1111111111000010100100,
    22'b0000000000001010001111,
    22'b0000000001011100001010,
    22'b0000000011001100110011,
    22'b0000000100101000111101,
    22'b0000000110000101001000,
    22'b0000000111010111000011,
    22'b0000001000110011001101,
    22'b0000001111100001010010,
    22'b0000010001111010111000,
    22'b0000010100011110101110,
    22'b0000011000001010001111,
    22'b0000011010011001100110,
    22'b0000011011001100110011,
    22'b0000011011010111000011,
    22'b0000011011101011100001,
    22'b0000011100011110101110,
    22'b0000011101000111101100,
    22'b0000011101111010111000,
    22'b0000011110000101001000,
    22'b0000011101110000101001,
    22'b0000011101010001111011,
    22'b0000011100101000111101,
    22'b0000011100001010001111,
    22'b0000011100001010001111,
    22'b0000011100110011001101,
    22'b0000011101100110011010,
    22'b0000011111000010100100,
    22'b0000100000010100011111,
    22'b0000100010000101001000,
    22'b0000100100001010001111,
    22'b0000100111000010100100,
    22'b0000101001010001111011,
    22'b0000101011101011100001,
    22'b0000101110000101001000,
    22'b0000110001011100001010,
    22'b0000110100000000000000,
    22'b0000110110001111010111,
    22'b0000111000010100011111,
    22'b0000111010000101001000,
    22'b0000111010111000010100,
    22'b0000111011010111000011,
    22'b0000111011100001010010,
    22'b0000111011101011100001,
    22'b0000111100010100011111,
    22'b0001000011100001010010,
    22'b0001000100101000111101,
    22'b0001000011110101110001,
    22'b0001000001110000101001,
    22'b0000111110101110000101,
    22'b0000111011001100110011,
    22'b0000110101110000101001,
    22'b0000110001110000101001,
    22'b0000101110011001100110,
    22'b0000101011110101110001,
    22'b0000101010000101001000,
    22'b0000101001011100001010,
    22'b0000101001011100001010,
    22'b0000101001100110011010,
    22'b0000101010100011110110,
    22'b0000101011100001010010,
    22'b0000101101000111101100,
    22'b0000101110101110000101,
    22'b0000110001011100001010,
    22'b0000110011100001010010,
    22'b0000110101110000101001,
    22'b0000110111110101110001,
    22'b0000111010001111010111,
    22'b0000111011100001010010,
    22'b0000111100001010001111,
    22'b0000111100110011001101,
    22'b0000111101100110011010,
    22'b0000111110011001100110,
    22'b0000111111101011100001,
    22'b0001000001000111101100,
    22'b0001000011101011100001,
    22'b0001000110011001100110,
    22'b0001001001011100001010,
    22'b0001001100111101011100,
    22'b0001010000101000111101,
    22'b0001010101100110011010,
    22'b0001011000111101011100,
    22'b0001011011100001010010,
    22'b0001011100101000111101,
    22'b0001010101100110011010,
    22'b0001010011010111000011,
    22'b0001010001010001111011,
    22'b0001001110100011110110,
    22'b0001001100101000111101,
    22'b0001001010111000010100,
    22'b0001001001100110011010,
    22'b0001000111110101110001,
    22'b0001000110100011110110,
    22'b0001000101011100001010,
    22'b0001000100001010001111,
    22'b0001000010100011110110,
    22'b0001000001010001111011,
    22'b0000111111110101110001,
    22'b0000111110000101001000,
    22'b0000111101010001111011,
    22'b0000111101000111101100,
    22'b0000111101100110011010,
    22'b0000111111010111000011,
    22'b0001000001011100001010,
    22'b0001000011110101110001,
    22'b0001000110100011110110,
    22'b0001001010000101001000,
    22'b0001001100011110101110,
    22'b0001001110111000010100,
    22'b0001010001000111101100,
    22'b0001010011101011100001,
    22'b0001010101011100001010,
    22'b0001010111001100110011,
    22'b0001011000101000111101,
    22'b0001011010100011110110,
    22'b0001011100000000000000,
    22'b0001011101100110011010,
    22'b0001011111100001010010,
    22'b0001100001111010111000,
    22'b0001100011001100110011,
    22'b0001100100000000000000,
    22'b0001100100101000111101,
    22'b0001100100011110101110,
    22'b0001100011110101110001,
    22'b0001100011000010100100,
    22'b0001100001100110011010,
    22'b0001011100000000000000,
    22'b0001011010011001100110,
    22'b0001011000010100011111,
    22'b0001010110101110000101,
    22'b0001010101010001111011,
    22'b0001010011101011100001,
    22'b0001010001111010111000,
    22'b0001010000111101011100,
    22'b0001010000010100011111,
    22'b0001010000001010001111,
    22'b0001010000101000111101,
    22'b0001010001010001111011,
    22'b0001010010000101001000,
    22'b0001010010111000010100,
    22'b0001010100000000000000,
    22'b0001010100110011001101,
    22'b0001010101011100001010,
    22'b0001010110001111010111,
    22'b0001010111100001010010,
    22'b0001011000011110101110,
    22'b0001011001100110011010,
    22'b0001011010111000010100,
    22'b0001011100000000000000,
    22'b0001011100011110101110,
    22'b0001011100101000111101,
    22'b0001011100101000111101,
    22'b0001011100110011001101,
    22'b0001011101000111101100,
    22'b0001011101111010111000,
    22'b0001011110111000010100,
    22'b0001100000010100011111,
    22'b0001100001010001111011,
    22'b0001100001111010111000,
    22'b0001100010011001100110,
    22'b0001100010101110000101,
    22'b0001100010111000010100,
    22'b0001100010111000010100,
    22'b0001100010101110000101,
    22'b0001100010001111010111,
    22'b0001100001011100001010,
    22'b0001100000011110101110,
    22'b0001011111000010100100,
    22'b0001011101000111101100,
    22'b0001011010011001100110,
    22'b0001011000011110101110,
    22'b0001010110100011110110,
    22'b0001010100110011001101,
    22'b0001010010111000010100,
    22'b0001010001010001111011,
    22'b0001010000000000000000,
    22'b0001001110100011110110,
    22'b0001001100011110101110,
    22'b0001001011101011100001,
    22'b0001001011010111000011,
    22'b0001001011100001010010,
    22'b0001001010111000010100,
    22'b0001001010111000010100,
    22'b0001001011000010100100,
    22'b0001001011101011100001,
    22'b0001001100010100011111,
    22'b0001001101011100001010,
    22'b0001001110111000010100,
    22'b0001001111110101110001,
    22'b0001010000010100011111,
    22'b0001010000101000111101,
    22'b0001010000110011001101,
    22'b0001010000110011001101,
    22'b0001010000010100011111,
    22'b0001001111101011100001,
    22'b0001001110111000010100,
    22'b0001001101111010111000,
    22'b0001001100101000111101,
    22'b0001001011110101110001,
    22'b0001001011100001010010,
    22'b0001001011101011100001,
    22'b0001001101011100001010,
    22'b0001001101000111101100,
    22'b0001001011100001010010,
    22'b0001001001100110011010,
    22'b0001000111101011100001,
    22'b0001000100110011001101,
    22'b0001000010100011110110,
    22'b0001000000010100011111,
    22'b0000111110011001100110,
    22'b0000111100011110101110,
    22'b0000111011110101110001,
    22'b0000111011110101110001,
    22'b0000111100010100011111,
    22'b0000111101000111101100,
    22'b0000111110101110000101,
    22'b0001000000011110101110,
    22'b0001000010101110000101,
    22'b0001000101010001111011,
    22'b0001001000110011001101,
    22'b0001001011101011100001,
    22'b0001001111000010100100,
    22'b0001010010101110000101,
    22'b0001010110101110000101,
    22'b0001011100000000000000,
    22'b0001011111101011100001,
    22'b0001100011001100110011,
    22'b0001100110100011110110,
    22'b0001101001110000101001,
    22'b0001101011110101110001,
    22'b0001101101010001111011,
    22'b0001101110001111010111,
    22'b0001101110100011110110,
    22'b0001101101111010111000,
    22'b0001101101010001111011,
    22'b0001101100001010001111,
    22'b0001101011001100110011,
    22'b0001101001010001111011,
    22'b0001100111110101110001,
    22'b0001100110101110000101,
    22'b0001100101111010111000,
    22'b0001100101011100001010,
    22'b0001100101000111101100,
    22'b0001100101010001111011,
    22'b0001100101011100001010,
    22'b0001100101011100001010,
    22'b0001100101100110011010,
    22'b0001100101100110011010,
    22'b0001100100101000111101,
    22'b0001100011101011100001,
    22'b0001100010011001100110,
    22'b0001100001000111101100,
    22'b0001011111101011100001,
    22'b0001011110100011110110,
    22'b0001011101100110011010,
    22'b0001011100011110101110,
    22'b0001011011010111000011,
    22'b0001011010011001100110,
    22'b0001011001011100001010,
    22'b0001011000010100011111,
    22'b0001010111110101110001,
    22'b0001010111010111000011,
    22'b0001010110011001100110,
    22'b0001010100111101011100,
    22'b0001010100001010001111,
    22'b0001010011101011100001,
    22'b0001010011100001010010,
    22'b0001010011110101110001,
    22'b0001010100010100011111,
    22'b0001010100011110101110,
    22'b0001010101000111101100,
    22'b0001010101111010111000,
    22'b0001010110111000010100,
    22'b0001010111000010100100,
    22'b0001010110111000010100,
    22'b0001010110011001100110,
    22'b0001010101100110011010,
    22'b0001010100010100011111,
    22'b0001010010101110000101,
    22'b0001010001000111101100,
    22'b0001001111010111000011,
    22'b0001001110101110000101,
    22'b0001001101110000101001,
    22'b0001001100110011001101,
    22'b0001001011010111000011,
    22'b0001001000010100011111,
    22'b0001000101011100001010,
    22'b0001000011001100110011,
    22'b0001000001011100001010,
    22'b0000111110011001100110,
    22'b0000111101110000101001,
    22'b0000111101000111101100,
    22'b0000111100000000000000,
    22'b0000111010101110000101,
    22'b0000111001100110011010,
    22'b0000110111101011100001,
    22'b0000110101110000101001,
    22'b0000110010111000010100,
    22'b0000110000110011001101,
    22'b0000101110100011110110,
    22'b0000101100101000111101,
    22'b0000101011010111000011,
    22'b0000101010111000010100,
    22'b0000101011010111000011,
    22'b0000101100010100011111,
    22'b0000101101100110011010,
    22'b0000101110111000010100,
    22'b0000110010101110000101,
    22'b0000110101010001111011,
    22'b0000110111100001010010,
    22'b0000111001111010111000,
    22'b0000111100000000000000,
    22'b0000111110011001100110,
    22'b0001000001010001111011,
    22'b0001000100110011001101,
    22'b0001001001110000101001,
    22'b0001001101010001111011,
    22'b0001010000001010001111,
    22'b0001010010111000010100,
    22'b0001010100110011001101,
    22'b0001010110100011110110,
    22'b0001010111001100110011,
    22'b0001010111010111000011,
    22'b0001010111010111000011,
    22'b0001010110101110000101,
    22'b0001010101011100001010,
    22'b0001010100011110101110,
    22'b0001010011001100110011,
    22'b0001010001011100001010,
    22'b0001001110100011110110,
    22'b0001001100010100011111,
    22'b0001001010011001100110,
    22'b0001001000110011001101,
    22'b0001000111100001010010,
    22'b0001000111101011100001,
    22'b0001001000001010001111,
    22'b0001001001000111101100,
    22'b0001001010000101001000,
    22'b0001001011101011100001,
    22'b0001001011110101110001,
    22'b0001001011100001010010,
    22'b0001001011000010100100,
    22'b0001001001100110011010,
    22'b0001001000000000000000,
    22'b0001000110100011110110,
    22'b0001000101010001111011,
    22'b0001000100101000111101,
    22'b0001000100011110101110,
    22'b0001000100011110101110,
    22'b0001000100011110101110,
    22'b0001000101000111101100,
    22'b0001000110001111010111,
    22'b0001000111101011100001,
    22'b0001001001010001111011,
    22'b0001001010000101001000,
    22'b0001001010100011110110,
    22'b0001001101011100001010,
    22'b0001001110101110000101,
    22'b0001001110101110000101,
    22'b0001001110000101001000,
    22'b0001001011000010100100,
    22'b0001000111110101110001,
    22'b0001000100000000000000,
    22'b0001000000001010001111,
    22'b0000111011100001010010,
    22'b0000110111000010100100,
    22'b0000110010001111010111,
    22'b0000101101100110011010,
    22'b0000100111110101110001,
    22'b0000011110000101001000,
    22'b0000010110100011110110,
    22'b0000010000011110101110,
    22'b0000001100000000000000,
    22'b0000000111110101110001,
    22'b0000000100110011001101,
    22'b0000000110000101001000,
    22'b0000001000011110101110,
    22'b0000001011110101110001,
    22'b0000001110011001100110,
    22'b0000010000101000111101,
    22'b0000010010011001100110,
    22'b0000010100011110101110,
    22'b0000010101100110011010,
    22'b0000010111000010100100,
    22'b0000010111110101110001,
    22'b0000011001100110011010,
    22'b0000011011101011100001,
    22'b0000011100010100011111,
    22'b0000011101111010111000,
    22'b0000011100011110101110,
    22'b0000011010001111010111,
    22'b0000011000001010001111,
    22'b0000010101010001111011,
    22'b0000010011000010100100,
    22'b0000010001110000101001,
    22'b0000010001010001111011,
    22'b0000010001011100001010,
    22'b0000010001111010111000,
    22'b0000010010011001100110,
    22'b0000010010001111010111,
    22'b0000010001111010111000,
    22'b0000010000001010001111,
    22'b0000001101010001111011,
    22'b0000001010101110000101,
    22'b0000000111000010100100,
    22'b0000000011110101110001,
    22'b1111111101100110011010,
    22'b1111111011010111000011,
    22'b1111110111110101110001,
    22'b1111110100111101011100,
    22'b1111110010111000010100,
    22'b1111110000111101011100,
    22'b1111101110111000010100,
    22'b1111100111010111000011,
    22'b1111100101100110011010,
    22'b1111100100111101011100,
    22'b1111100100001010001111,
    22'b1111100010101110000101,
    22'b1111100001011100001010,
    22'b1111100000000000000000,
    22'b1111011101010001111011,
    22'b1111011100110011001101,
    22'b1111011011000010100100,
    22'b1111011001000111101100,
    22'b1111010111000010100100,
    22'b1111010111001100110011,
    22'b1111010111110101110001,
    22'b1111011000001010001111,
    22'b1111010111010111000011,
    22'b1111011000101000111101,
    22'b1111011001110000101001,
    22'b1111011010001111010111,
    22'b1111011011000010100100,
    22'b1111011100000000000000,
    22'b1111011100111101011100,
    22'b1111011101000111101100,
    22'b1111011101011100001010,
    22'b1111011100101000111101,
    22'b1111011011010111000011,
    22'b1111011001010001111011,
    22'b1111010111010111000011,
    22'b1111010100111101011100,
    22'b1111001010011001100110,
    22'b1111000100001010001111,
    22'b1111000000110011001101,
    22'b1110111010000101001000,
    22'b1110110011000010100100,
    22'b1110110001100110011010,
    22'b1110110000001010001111,
    22'b1110110000011110101110,
    22'b1110110100001010001111,
    22'b1110110101111010111000,
    22'b1110110111001100110011,
    22'b1110111000000000000000,
    22'b1110111001000111101100,
    22'b1110111010001111010111,
    22'b1110111100001010001111,
    22'b1110111110111000010100,
    22'b1111000011001100110011,
    22'b1111000110101110000101,
    22'b1111001001110000101001,
    22'b1111001101110000101001,
    22'b1111010001010001111011,
    22'b1111010100110011001101,
    22'b1111011000011110101110,
    22'b1111011101011100001010,
    22'b1111100001000111101100,
    22'b1111100100101000111101,
    22'b1111101110111000010100,
    22'b1111101111001100110011,
    22'b1111101110111000010100,
    22'b1111101100110011001101,
    22'b1111101010011001100110,
    22'b1111101000001010001111,
    22'b1111100101000111101100,
    22'b1111100001010001111011,
    22'b1111011111000010100100,
    22'b1111011101000111101100,
    22'b1111011011101011100001,
    22'b1111011011010111000011,
    22'b1111011011101011100001,
    22'b1111011011110101110001,
    22'b1111011110001111010111,
    22'b1111100000000000000000,
    22'b1111100001111010111000,
    22'b1111100011101011100001,
    22'b1111100100101000111101,
    22'b1111100100101000111101,
    22'b1111100101011100001010,
    22'b1111100110111000010100,
    22'b1111100111101011100001,
    22'b1111101000111101011100,
    22'b1111101010000101001000,
    22'b1111101011001100110011,
    22'b1111101011101011100001,
    22'b1111101011101011100001,
    22'b1111101011000010100100,
    22'b1111101001111010111000,
    22'b1111100100110011001101,
    22'b1111100010111000010100,
    22'b1111100000011110101110,
    22'b1111011110111000010100,
    22'b1111011101100110011010,
    22'b1111011100000000000000,
    22'b1111011010101110000101,
    22'b1111011001100110011010,
    22'b1111011000010100011111,
    22'b1111010110101110000101,
    22'b1111010101111010111000,
    22'b1111010101110000101001,
    22'b1111010101111010111000,
    22'b1111010110101110000101,
    22'b1111010111001100110011,
    22'b1111010111110101110001,
    22'b1111011000001010001111,
    22'b1111011000001010001111,
    22'b1111011000001010001111,
    22'b1111010111110101110001,
    22'b1111010111100001010010,
    22'b1111010111000010100100,
    22'b1111010111000010100100,
    22'b1111010110111000010100,
    22'b1111010110101110000101,
    22'b1111010110000101001000,
    22'b1111010100111101011100,
    22'b1111010011001100110011,
    22'b1111001111110101110001,
    22'b1111001100011110101110,
    22'b1111001000111101011100,
    22'b1111000100110011001101,
    22'b1110111110100011110110,
    22'b1110111001111010111000,
    22'b1110110101110000101001,
    22'b1110100100110011001101,
    22'b1110100011001100110011,
    22'b1110100011001100110011,
    22'b1110100101010001111011,
    22'b1110100111010111000011,
    22'b1110101010001111010111,
    22'b1110101101111010111000,
    22'b1110110011100001010010,
    22'b1110110111100001010010,
    22'b1110111010111000010100,
    22'b1110111101110000101001,
    22'b1111000001100110011010,
    22'b1111000011110101110001,
    22'b1111000110001111010111,
    22'b1111001000010100011111,
    22'b1111001011000010100100,
    22'b1111001101000111101100,
    22'b1111001111001100110011,
    22'b1111010001010001111011,
    22'b1111010011101011100001,
    22'b1111010101100110011010,
    22'b1111010111100001010010,
    22'b1111011001110000101001,
    22'b1111011010111000010100,
    22'b1111011011110101110001,
    22'b1111011100101000111101,
    22'b1111011101011100001010,
    22'b1111011101111010111000,
    22'b1111011110001111010111,
    22'b1111011110101110000101,
    22'b1111011111001100110011,
    22'b1111011111101011100001,
    22'b1111100000011110101110,
    22'b1111100001010001111011,
    22'b1111100010011001100110,
    22'b1111100011001100110011,
    22'b1111100011110101110001,
    22'b1111100011101011100001,
    22'b1111100010011001100110,
    22'b1111100000111101011100,
    22'b1111100000011110101110,
    22'b1111100001000111101100,
    22'b1111101001000111101100,
    22'b1111101010000101001000,
    22'b1111101010001111010111,
    22'b1111101001111010111000,
    22'b1111101010100011110110,
    22'b1111101101110000101001,
    22'b1111101111101011100001,
    22'b1111110001100110011010,
    22'b1111110001111010111000,
    22'b1111110100111101011100,
    22'b1111111010000101001000,
    22'b1111111101000111101100,
    22'b0000000000011110101110,
    22'b0000000001111010111000,
    22'b0000000010000101001000,
    22'b0000000010101110000101,
    22'b0000000100010100011111,
    22'b0000000101010001111011,
    22'b0000000100110011001101,
    22'b0000000101100110011010,
    22'b0000000110000101001000,
    22'b0000000101010001111011,
    22'b0000000101010001111011,
    22'b0000000100111101011100,
    22'b0000000011110101110001,
    22'b0000000001000111101100,
    22'b1111111100110011001101,
    22'b1111111010001111010111,
    22'b1111110111110101110001,
    22'b1111110110001111010111,
    22'b1111110101111010111000,
    22'b1111110100010100011111,
    22'b1111110010000101001000,
    22'b1111101101110000101001,
    22'b1111101000111101011100,
    22'b1111100011100001010010,
    22'b1111011110000101001000,
    22'b1111011011000010100100,
    22'b1111011100011110101110,
    22'b1111100000011110101110,
    22'b1111100010011001100110,
    22'b1111100100001010001111,
    22'b1111100110101110000101,
    22'b1111100111010111000011,
    22'b1111101000010100011111,
    22'b1111101001000111101100,
    22'b1111101001111010111000,
    22'b1111101011100001010010,
    22'b1111101100101000111101,
    22'b1111101101000111101100,
    22'b1111101101111010111000,
    22'b1111101110001111010111,
    22'b1111101110111000010100,
    22'b1111101111110101110001,
    22'b1111110000111101011100,
    22'b1111110001000111101100,
    22'b1111110000101000111101,
    22'b1111110001000111101100,
    22'b1111110000001010001111,
    22'b1111101110100011110110,
    22'b1111101011110101110001,
    22'b1111101001110000101001,
    22'b1111100110101110000101,
    22'b1111100101010001111011,
    22'b1111100011000010100100,
    22'b1111100010000101001000,
    22'b1111100000111101011100,
    22'b1111011111110101110001,
    22'b1111100001010001111011,
    22'b1111100001000111101100,
    22'b1111011111110101110001,
    22'b1111100010111000010100,
    22'b1111100000010100011111,
    22'b1111001110000101001000,
    22'b1111010100000000000000,
    22'b1111011010101110000101,
    22'b1111100001100110011010,
    22'b1111100110000101001000,
    22'b1111101001111010111000,
    22'b1111101101000111101100,
    22'b1111110000111101011100,
    22'b1111110010100011110110,
    22'b1111110011110101110001,
    22'b1111110100110011001101,
    22'b1111110110000101001000,
    22'b1111110111010111000011,
    22'b1111111000010100011111,
    22'b1111111001011100001010,
    22'b1111111010011001100110,
    22'b1111111010101110000101,
    22'b1111111010111000010100,
    22'b1111111010011001100110,
    22'b1111111010100011110110,
    22'b1111111001110000101001,
    22'b1111111000111101011100,
    22'b1111110111010111000011,
    22'b1111110110001111010111,
    22'b1111110101011100001010,
    22'b1111110101011100001010,
    22'b1111110110111000010100,
    22'b1111110110011001100110,
    22'b1111111000101000111101,
    22'b1111111000101000111101,
    22'b1111110110101110000101,
    22'b1111110011000010100100,
    22'b1111101110111000010100,
    22'b1111101001011100001010,
    22'b1111101101110000101001,
    22'b1111101111000010100100,
    22'b1111110000001010001111,
    22'b1111110011010111000011,
    22'b1111110011101011100001,
    22'b1111110000010100011111,
    22'b1111101101111010111000,
    22'b1111101101100110011010,
    22'b1111110010011001100110,
    22'b1111110000111101011100,
    22'b1111101111001100110011,
    22'b1111110010000101001000,
    22'b1111110011110101110001,
    22'b1111110011101011100001,
    22'b1111110011000010100100,
    22'b1111110001010001111011,
    22'b1111110000011110101110,
    22'b1111110001110000101001,
    22'b1111101101000111101100,
    22'b1111100011110101110001,
    22'b1111010111001100110011,
    22'b1111000110111000010100,
    22'b1110111011100001010010,
    22'b1110101100110011001101,
    22'b1110011001011100001010,
    22'b1110001111101011100001,
    22'b1110000110000101001000,
    22'b1101111101111010111000,
    22'b1101111000000000000000,
    22'b1101110111100001010010,
    22'b1101111000101000111101,
    22'b1101111100010100011111,
    22'b1110000010011001100110,
    22'b1110001000101000111101,
    22'b1110001110101110000101,
    22'b1110010111000010100100,
    22'b1110100101010001111011,
    22'b1110100111010111000011,
    22'b1110101011000010100100,
    22'b1110101110000101001000,
    22'b1110110001000111101100,
    22'b1110110100000000000000,
    22'b1110110110101110000101,
    22'b1110111000001010001111,
    22'b1110111000111101011100,
    22'b1110111000111101011100,
    22'b1110111000000000000000,
    22'b1110110110101110000101,
    22'b1110110101000111101100,
    22'b1110110011001100110011,
    22'b1110110010000101001000,
    22'b1110110001000111101100,
    22'b1110110000011110101110,
    22'b1110110000001010001111,
    22'b1110110000001010001111,
    22'b1110110000101000111101,
    22'b1110110001110000101001,
    22'b1110110010101110000101,
    22'b1110110100000000000000,
    22'b1110110101010001111011,
    22'b1110110111100001010010,
    22'b1110111001010001111011,
    22'b1110111010111000010100,
    22'b1110111100011110101110,
    22'b1110111110011001100110,
    22'b1110111111100001010010,
    22'b1111000000101000111101,
    22'b1111000001110000101001,
    22'b1111000001111010111000,
    22'b1111000001011100001010,
    22'b1111000000101000111101,
    22'b1111000000000000000000,
    22'b1110111111101011100001,
    22'b1110111111010111000011,
    22'b1110111111000010100100,
    22'b1110111110100011110110,
    22'b1110111110000101001000,
    22'b1110111101010001111011,
    22'b1110111100001010001111,
    22'b1110111010111000010100,
    22'b1110111001010001111011,
    22'b1110110111010111000011,
    22'b1110110101110000101001,
    22'b1110110100000000000000,
    22'b1110110010001111010111,
    22'b1110110000001010001111,
    22'b1110101111000010100100,
    22'b1110101110001111010111,
    22'b1110101101011100001010,
    22'b1110101100111101011100,
    22'b1110101100110011001101,
    22'b1110101100010100011111,
    22'b1110101100111101011100,
    22'b1110101100101000111101,
    22'b1110101011101011100001,
    22'b1110101011100001010010,
    22'b1110101101100110011010,
    22'b1110101111000010100100,
    22'b1110110000111101011100,
    22'b1110111110111000010100,
    22'b1111000001011100001010,
    22'b1111000011101011100001,
    22'b1111000101110000101001,
    22'b1111001000000000000000,
    22'b1111001001000111101100,
    22'b1111001001111010111000,
    22'b1111001010100011110110,
    22'b1111001011001100110011,
    22'b1111001010011001100110,
    22'b1111001000111101011100,
    22'b1111000110100011110110,
    22'b1111000100111101011100,
    22'b1111000011100001010010,
    22'b1111000010001111010111,
    22'b1110111111110101110001,
    22'b1110111101011100001010,
    22'b1110111011000010100100,
    22'b1110110111010111000011,
    22'b1110110100001010001111,
    22'b1110110001000111101100,
    22'b1110101111001100110011,
    22'b1110101101011100001010,
    22'b1110101011010111000011,
    22'b1110101001110000101001,
    22'b1110101000110011001101,
    22'b1110101000010100011111,
    22'b1110101000011110101110,
    22'b1110101001011100001010,
    22'b1110101010100011110110,
    22'b1110101011000010100100,
    22'b1110101110001111010111,
    22'b1110110001011100001010,
    22'b1110110100000000000000,
    22'b1110110110111000010100,
    22'b1110111001011100001010,
    22'b1110111100011110101110,
    22'b1110111110101110000101,
    22'b1111000001000111101100,
    22'b1111000100010100011111,
    22'b1111000110000101001000,
    22'b1111000111010111000011,
    22'b1111000111100001010010,
    22'b1111000110101110000101,
    22'b1111000101010001111011,
    22'b1111000011100001010010,
    22'b1111000001110000101001,
    22'b1110111111001100110011,
    22'b1110111101011100001010,
    22'b1110111100011110101110,
    22'b1110111100011110101110,
    22'b1110111101111010111000,
    22'b1110111111110101110001,
    22'b1111000001111010111000,
    22'b1111000100011110101110,
    22'b1111001001110000101001,
    22'b1111001010111000010100,
    22'b1111001100001010001111,
    22'b1111001100111101011100,
    22'b1111001110000101001000,
    22'b1111001111001100110011,
    22'b1111010000111101011100,
    22'b1111010010100011110110,
    22'b1111010100001010001111,
    22'b1111010101011100001010,
    22'b1111010101100110011010,
    22'b1111010101010001111011,
    22'b1111010100101000111101,
    22'b1111010100001010001111,
    22'b1111010100001010001111,
    22'b1111010011110101110001,
    22'b1111010010111000010100,
    22'b1111010001000111101100,
    22'b1111010000000000000000,
    22'b1111001111100001010010,
    22'b1111001111100001010010,
    22'b1111001111100001010010,
    22'b1111001111010111000011,
    22'b1111001111110101110001,
    22'b1111010001100110011010,
    22'b1111011001010001111011,
    22'b1111011010101110000101,
    22'b1111011100111101011100,
    22'b1111011111000010100100,
    22'b1111100001000111101100,
    22'b1111100010111000010100,
    22'b1111100101010001111011,
    22'b1111100111010111000011,
    22'b1111101001010001111011,
    22'b1111101011000010100100,
    22'b1111101100111101011100,
    22'b1111101110011001100110,
    22'b1111110000010100011111,
    22'b1111110010011001100110,
    22'b1111110101000111101100,
    22'b1111110111100001010010,
    22'b1111111010011001100110,
    22'b1111111101110000101001,
    22'b0000000011101011100001,
    22'b0000000111000010100100,
    22'b0000001001000111101100,
    22'b0000001011010111000011,
    22'b0000001101110000101001,
    22'b0000001111010111000011,
    22'b0000010000110011001101,
    22'b0000010010100011110110,
    22'b0000010100011110101110,
    22'b0000010101011100001010,
    22'b0000010101110000101001,
    22'b0000010101100110011010,
    22'b0000010100111101011100,
    22'b0000010100101000111101,
    22'b0000010000101000111101,
    22'b0000010010000101001000,
    22'b0000010100010100011111,
    22'b0000010111001100110011,
    22'b0000011001111010111000,
    22'b0000011101000111101100,
    22'b0000011110111000010100,
    22'b0000011111110101110001,
    22'b0000100000011110101110,
    22'b0000100000111101011100,
    22'b0000100001011100001010,
    22'b0000100001111010111000,
    22'b0000100010111000010100,
    22'b0000100100101000111101,
    22'b0000100110000101001000,
    22'b0000100111110101110001,
    22'b0000101001110000101001,
    22'b0000101100001010001111,
    22'b0000101101100110011010,
    22'b0000101111000010100100,
    22'b0000101111101011100001,
    22'b0000101111010111000011,
    22'b0000101111101011100001,
    22'b0000110000000000000000,
    22'b0000110000000000000000,
    22'b0000110000101000111101,
    22'b0000110010011001100110,
    22'b0000110011101011100001,
    22'b0000110011000010100100,
    22'b0000110100010100011111,
    22'b0000110011101011100001,
    22'b0000011001100110011010,
    22'b0000001000001010001111,
    22'b1111111000010100011111,
    22'b1111101001000111101100,
    22'b1111011010101110000101,
    22'b1111010011110101110001,
    22'b1111010000111101011100,
    22'b1111010000110011001101,
    22'b1111010101010001111011,
    22'b1111011010111000010100,
    22'b1111100000101000111101,
    22'b1111101000010100011111,
    22'b1111101101000111101100,
    22'b1111110000110011001101,
    22'b1111110011001100110011,
    22'b1111110100110011001101,
    22'b1111110101011100001010,
    22'b1111110101110000101001,
    22'b1111110110011001100110,
    22'b1111110110100011110110,
    22'b1111110110101110000101,
    22'b1111110110111000010100,
    22'b1111110111010111000011,
    22'b1111111011100001010010,
    22'b1111111101010001111011,
    22'b0000000000001010001111,
    22'b0000000010101110000101,
    22'b0000000101100110011010,
    22'b0000001000011110101110,
    22'b0000001100110011001101,
    22'b0000010000001010001111,
    22'b0000010011010111000011,
    22'b0000010100111101011100,
    22'b0000011000011110101110,
    22'b0000011011001100110011,
    22'b0000011110011001100110,
    22'b0000100001110000101001,
    22'b0000100111001100110011,
    22'b0000101011101011100001,
    22'b0000101111000010100100,
    22'b0000110011110101110001,
    22'b0000110110011001100110,
    22'b0000110110101110000101,
    22'b0000110110001111010111,
    22'b0000110011010111000011,
    22'b0000110000000000000000,
    22'b0000101011100001010010,
    22'b0000100110100011110110,
    22'b0000011111010111000011,
    22'b0000011010100011110110,
    22'b0000001100101000111101,
    22'b0000001010100011110110,
    22'b0000001001100110011010,
    22'b0000001010000101001000,
    22'b0000001011001100110011,
    22'b0000001100010100011111,
    22'b0000001100111101011100,
    22'b0000001101011100001010,
    22'b0000001101000111101100,
    22'b0000001110100011110110,
    22'b0000010000000000000000,
    22'b0000001111101011100001,
    22'b0000010001100110011010,
    22'b0000010100000000000000,
    22'b0000011000011110101110,
    22'b0000011101111010111000,
    22'b0000100010011001100110,
    22'b0000100111101011100001,
    22'b0000101100000000000000,
    22'b0000101111010111000011,
    22'b0000110100010100011111,
    22'b0000110111101011100001,
    22'b0000111010100011110110,
    22'b0000111100111101011100,
    22'b0001000000000000000000,
    22'b0001000010000101001000,
    22'b0001000010111000010100,
    22'b0001000011100001010010,
    22'b0001000100010100011111,
    22'b0001000100111101011100,
    22'b0001000100110011001101,
    22'b0001000100011110101110,
    22'b0001000100010100011111,
    22'b0001000011101011100001,
    22'b0000111110001111010111,
    22'b0000111100101000111101,
    22'b0000111011110101110001,
    22'b0000111011110101110001,
    22'b0000111011110101110001,
    22'b0000111010011001100110,
    22'b0000111000111101011100,
    22'b0000110111010111000011,
    22'b0000110100011110101110,
    22'b0000110001110000101001,
    22'b0000101110001111010111,
    22'b0000101001110000101001,
    22'b0000100011000010100100,
    22'b0000011101111010111000,
    22'b0000011000110011001101,
    22'b0000010100001010001111,
    22'b0000001110101110000101,
    22'b0000001011100001010010,
    22'b0000001001000111101100,
    22'b0000001000000000000000,
    22'b0000001000011110101110,
    22'b0000001010011001100110,
    22'b0000001100111101011100,
    22'b0000010000111101011100,
    22'b0000010100000000000000,
    22'b0000010111100001010010,
    22'b0000011011000010100100,
    22'b0000011111000010100100,
    22'b0000100001100110011010,
    22'b0000100011101011100001,
    22'b0000100101010001111011,
    22'b0000100111010111000011,
    22'b0000101000110011001101,
    22'b0000101010001111010111,
    22'b0000101011101011100001,
    22'b0000101100110011001101,
    22'b0000101101010001111011,
    22'b0000101101010001111011,
    22'b0000101011110101110001,
    22'b0000101010111000010100,
    22'b0000101000111101011100,
    22'b0000100110100011110110,
    22'b0000100011101011100001,
    22'b0000100001111010111000,
    22'b0000100000101000111101,
    22'b0000011111010111000011,
    22'b0000011101110000101001,
    22'b0000011100101000111101,
    22'b0000011100000000000000,
    22'b0000011011110101110001,
    22'b0000011100111101011100,
    22'b0000011110001111010111,
    22'b0000011111100001010010,
    22'b0000100000010100011111,
    22'b0000100000111101011100,
    22'b0000100001010001111011,
    22'b0000100001010001111011,
    22'b0000100000110011001101,
    22'b0000100000000000000000,
    22'b0000011111010111000011,
    22'b0000011111000010100100,
    22'b0000011111010111000011,
    22'b0000011111101011100001,
    22'b0000100000000000000000,
    22'b0000100000101000111101,
    22'b0000100001110000101001,
    22'b0000100011001100110011,
    22'b0000100101011100001010,
    22'b0000101000000000000000,
    22'b0000101100101000111101,
    22'b0000110000010100011111,
    22'b0000110011101011100001,
    22'b0000110110100011110110,
    22'b0000111000110011001101,
    22'b0000111001100110011010,
    22'b0000111010000101001000,
    22'b0000111010100011110110,
    22'b0000111011101011100001,
    22'b0000111100111101011100,
    22'b0000111110111000010100,
    22'b0001001011001100110011,
    22'b0001001100110011001101,
    22'b0001001101110000101001,
    22'b0001010000000000000000,
    22'b0001010001110000101001,
    22'b0001010011010111000011,
    22'b0001010100101000111101,
    22'b0001010110000101001000,
    22'b0001011000001010001111,
    22'b0001011001010001111011,
    22'b0001011001111010111000,
    22'b0001011011000010100100,
    22'b0001011101100110011010,
    22'b0001011110001111010111,
    22'b0001011111000010100100,
    22'b0001100000111101011100,
    22'b0001100001100110011010,
    22'b0001100001111010111000,
    22'b0001100010000101001000,
    22'b0001100001100110011010,
    22'b0001011110101110000101,
    22'b0001011100010100011111,
    22'b0001011001110000101001,
    22'b0001010111100001010010,
    22'b0001010100101000111101,
    22'b0001010010101110000101,
    22'b0001010001000111101100,
    22'b0001001111100001010010,
    22'b0001001101010001111011,
    22'b0001001011100001010010,
    22'b0001001001011100001010,
    22'b0001000111000010100100,
    22'b0001000100011110101110,
    22'b0001000010101110000101,
    22'b0001000001011100001010,
    22'b0001000000011110101110,
    22'b0000111111110101110001,
    22'b0000111111000010100100,
    22'b0000111110100011110110,
    22'b0000111110011001100110,
    22'b0000111110011001100110,
    22'b0000111111001100110011,
    22'b0000111111110101110001,
    22'b0001000000001010001111,
    22'b0001000000010100011111,
    22'b0001000000001010001111,
    22'b0001000000010100011111,
    22'b0001000001000111101100,
    22'b0001000010001111010111,
    22'b0001000100001010001111,
    22'b0001000110111000010100,
    22'b0001001000111101011100,
    22'b0001001011010111000011,
    22'b0001001101111010111000,
    22'b0001010000111101011100,
    22'b0001010011001100110011,
    22'b0001010101100110011010,
    22'b0001010111001100110011,
    22'b0001011000001010001111,
    22'b0001011001100110011010,
    22'b0001011010011001100110,
    22'b0001011010101110000101,
    22'b0001011011001100110011,
    22'b0001011011100001010010,
    22'b0001011011001100110011,
    22'b0001011010100011110110
};

parameter logic signed [`GYRO_WIDTH-1:0] WY_TEST_VECTOR[`NUM_ELEMENTS] = {
    22'b0000000101110000101001,
    22'b0000000101000111101100,
    22'b0000000100110011001101,
    22'b0000000100011110101110,
    22'b0000000100001010001111,
    22'b0000000011110101110001,
    22'b0000000011100001010010,
    22'b0000000011010111000011,
    22'b0000000011001100110011,
    22'b0000000010111000010100,
    22'b0000000010100011110110,
    22'b0000000010001111010111,
    22'b0000000001110000101001,
    22'b0000000001000111101100,
    22'b0000000000101000111101,
    22'b0000000000001010001111,
    22'b1111111111100001010010,
    22'b1111111110111000010100,
    22'b1111111110011001100110,
    22'b1111111101111010111000,
    22'b1111111101011100001010,
    22'b1111111100111101011100,
    22'b1111111100011110101110,
    22'b1111111100001010001111,
    22'b1111111011110101110001,
    22'b1111111011101011100001,
    22'b1111111011110101110001,
    22'b1111111100000000000000,
    22'b1111111100001010001111,
    22'b1111111100011110101110,
    22'b1111111100110011001101,
    22'b1111111101000111101100,
    22'b1111111101011100001010,
    22'b1111111101110000101001,
    22'b1111111110001111010111,
    22'b1111111110100011110110,
    22'b1111111110111000010100,
    22'b1111111111010111000011,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111101011100001,
    22'b1111111111010111000011,
    22'b1111111110101110000101,
    22'b1111111110000101001000,
    22'b1111111101011100001010,
    22'b1111111100111101011100,
    22'b1111111100101000111101,
    22'b1111111100011110101110,
    22'b1111111100011110101110,
    22'b1111111100101000111101,
    22'b1111111100111101011100,
    22'b1111111101010001111011,
    22'b1111111101110000101001,
    22'b1111111110000101001000,
    22'b1111111110011001100110,
    22'b1111111110111000010100,
    22'b1111111111010111000011,
    22'b1111111111101011100001,
    22'b1111111111110101110001,
    22'b0000000000001010001111,
    22'b0000000000010100011111,
    22'b0000000000101000111101,
    22'b0000000000110011001101,
    22'b0000000000110011001101,
    22'b0000000000001010001111,
    22'b1111111111001100110011,
    22'b1111111110111000010100,
    22'b1111111110011001100110,
    22'b1111111110000101001000,
    22'b1111111110001111010111,
    22'b1111111110111000010100,
    22'b1111111111100001010010,
    22'b0000000000001010001111,
    22'b0000000000011110101110,
    22'b0000000000101000111101,
    22'b0000000001011100001010,
    22'b0000000011110101110001,
    22'b0000000111100001010010,
    22'b0000001011010111000011,
    22'b0000010000111101011100,
    22'b0000011001111010111000,
    22'b0000011110101110000101,
    22'b0000100000011110101110,
    22'b0000100000010100011111,
    22'b0000011011101011100001,
    22'b0000010011100001010010,
    22'b0000001100101000111101,
    22'b0000000101111010111000,
    22'b0000000000001010001111,
    22'b1111111011000010100100,
    22'b1111111001010001111011,
    22'b1111111001110000101001,
    22'b1111111100000000000000,
    22'b1111111111110101110001,
    22'b0000000010111000010100,
    22'b0000000101011100001010,
    22'b0000000111101011100001,
    22'b0000001001011100001010,
    22'b0000001010001111010111,
    22'b0000001010100011110110,
    22'b0000001010001111010111,
    22'b0000001001010001111011,
    22'b0000000111100001010010,
    22'b0000000110101110000101,
    22'b0000000110000101001000,
    22'b0000000101010001111011,
    22'b0000000100001010001111,
    22'b0000000011101011100001,
    22'b0000000010100011110110,
    22'b0000000001111010111000,
    22'b0000000001011100001010,
    22'b0000000000110011001101,
    22'b0000000000101000111101,
    22'b0000000001000111101100,
    22'b0000000001100110011010,
    22'b0000000010001111010111,
    22'b0000000010011001100110,
    22'b0000000010100011110110,
    22'b0000000010011001100110,
    22'b0000000001111010111000,
    22'b0000000001010001111011,
    22'b0000000000110011001101,
    22'b0000000000001010001111,
    22'b1111111110101110000101,
    22'b1111111110001111010111,
    22'b1111111110101110000101,
    22'b1111111111000010100100,
    22'b1111111111000010100100,
    22'b1111111110101110000101,
    22'b1111111110100011110110,
    22'b1111111110001111010111,
    22'b1111111110000101001000,
    22'b1111111101100110011010,
    22'b1111111101010001111011,
    22'b1111111100101000111101,
    22'b1111111100001010001111,
    22'b1111111011010111000011,
    22'b1111111011010111000011,
    22'b1111111100000000000000,
    22'b1111111100101000111101,
    22'b1111111110001111010111,
    22'b0000000000000000000000,
    22'b0000000001011100001010,
    22'b0000000010001111010111,
    22'b0000000011000010100100,
    22'b0000000011010111000011,
    22'b0000000011110101110001,
    22'b0000000100010100011111,
    22'b0000000100011110101110,
    22'b0000000011000010100100,
    22'b0000000000110011001101,
    22'b1111111110100011110110,
    22'b1111111101000111101100,
    22'b1111111010011001100110,
    22'b1111111010000101001000,
    22'b1111111001010001111011,
    22'b1111111001100110011010,
    22'b1111111010000101001000,
    22'b1111111010011001100110,
    22'b1111111010101110000101,
    22'b1111111010111000010100,
    22'b1111111011001100110011,
    22'b1111111011110101110001,
    22'b1111111101000111101100,
    22'b1111111101111010111000,
    22'b1111111110001111010111,
    22'b1111111110100011110110,
    22'b1111111110000101001000,
    22'b1111111101110000101001,
    22'b1111111110000101001000,
    22'b1111111110101110000101,
    22'b1111111111001100110011,
    22'b0000000000000000000000,
    22'b0000000000011110101110,
    22'b0000000000101000111101,
    22'b0000000000110011001101,
    22'b1111111001011100001010,
    22'b1111110100000000000000,
    22'b1111110001000111101100,
    22'b1111101111001100110011,
    22'b1111101111010111000011,
    22'b1111101111001100110011,
    22'b1111101111100001010010,
    22'b1111110010000101001000,
    22'b1111101110000101001000,
    22'b1111101100101000111101,
    22'b1111101110000101001000,
    22'b1111110000011110101110,
    22'b1111111010000101001000,
    22'b0000000100000000000000,
    22'b0000001100110011001101,
    22'b0000010011010111000011,
    22'b0000011001010001111011,
    22'b0000011100001010001111,
    22'b0000011101110000101001,
    22'b0000011110101110000101,
    22'b0000011110101110000101,
    22'b0000011110111000010100,
    22'b0000011110001111010111,
    22'b0000011101111010111000,
    22'b0000011100000000000000,
    22'b0000010111101011100001,
    22'b0000010100000000000000,
    22'b0000010010111000010100,
    22'b0000010000011110101110,
    22'b0000001110101110000101,
    22'b0000010000110011001101,
    22'b0000010100110011001101,
    22'b0000011001100110011010,
    22'b0000011110000101001000,
    22'b0000100010111000010100,
    22'b0000100111001100110011,
    22'b0000101011001100110011,
    22'b0000110000011110101110,
    22'b0000110100000000000000,
    22'b0000110110001111010111,
    22'b0000110111100001010010,
    22'b0000110111101011100001,
    22'b0000110110100011110110,
    22'b0000110100010100011111,
    22'b0000110001000111101100,
    22'b0000101011001100110011,
    22'b0000100101011100001010,
    22'b0000011110101110000101,
    22'b0000010111001100110011,
    22'b0000001111101011100001,
    22'b0000000110000101001000,
    22'b1111111111100001010010,
    22'b1111111001110000101001,
    22'b1111110100101000111101,
    22'b1111101111000010100100,
    22'b1111101011101011100001,
    22'b1111101001010001111011,
    22'b1111100111110101110001,
    22'b1111100111001100110011,
    22'b1111100111101011100001,
    22'b1111101001000111101100,
    22'b1111101100010100011111,
    22'b1111101111100001010010,
    22'b1111110011000010100100,
    22'b1111110111000010100100,
    22'b1111111100010100011111,
    22'b0000000000010100011111,
    22'b0000000100001010001111,
    22'b0000000111001100110011,
    22'b0000001000010100011111,
    22'b0000001001100110011010,
    22'b0000001010011001100110,
    22'b0000000101110000101001,
    22'b1111111100101000111101,
    22'b1111111110101110000101,
    22'b1111111101111010111000,
    22'b1111111010111000010100,
    22'b1111110011110101110001,
    22'b1111101010000101001000,
    22'b1111100111000010100100,
    22'b1111100110001111010111,
    22'b1111101000110011001101,
    22'b1111101101000111101100,
    22'b1111101110111000010100,
    22'b1111101110100011110110,
    22'b1111101111110101110001,
    22'b1111110011000010100100,
    22'b1111110110101110000101,
    22'b1111111011101011100001,
    22'b0000000000010100011111,
    22'b0000000011110101110001,
    22'b0000000011110101110001,
    22'b0000000011010111000011,
    22'b0000000001100110011010,
    22'b0000000000111101011100,
    22'b0000000000110011001101,
    22'b1111111111100001010010,
    22'b1111111110001111010111,
    22'b1111111100010100011111,
    22'b1111111001011100001010,
    22'b1111110111110101110001,
    22'b1111110111001100110011,
    22'b1111110110111000010100,
    22'b1111110111100001010010,
    22'b1111111000001010001111,
    22'b1111111000111101011100,
    22'b1111111001111010111000,
    22'b1111111100000000000000,
    22'b1111111101110000101001,
    22'b1111111111100001010010,
    22'b0000000001011100001010,
    22'b0000000011000010100100,
    22'b0000000011100001010010,
    22'b0000000011110101110001,
    22'b0000000011110101110001,
    22'b0000000011101011100001,
    22'b0000000011001100110011,
    22'b0000000010100011110110,
    22'b0000000001100110011010,
    22'b0000000000010100011111,
    22'b1111111110011001100110,
    22'b1111111101010001111011,
    22'b1111111100010100011111,
    22'b1111111011101011100001,
    22'b1111111011001100110011,
    22'b1111111011000010100100,
    22'b1111111010111000010100,
    22'b1111111011000010100100,
    22'b1111111011101011100001,
    22'b1111111100010100011111,
    22'b1111111101010001111011,
    22'b1111111110000101001000,
    22'b1111111111001100110011,
    22'b1111111111110101110001,
    22'b0000000000011110101110,
    22'b0000000000110011001101,
    22'b0000000001010001111011,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001000111101100,
    22'b0000000000101000111101,
    22'b0000000000000000000000,
    22'b1111111111010111000011,
    22'b1111111110111000010100,
    22'b1111111110011001100110,
    22'b1111111101110000101001,
    22'b1111111101010001111011,
    22'b1111111101000111101100,
    22'b1111111100111101011100,
    22'b1111111100111101011100,
    22'b1111111101000111101100,
    22'b1111111101010001111011,
    22'b1111111101110000101001,
    22'b1111111110001111010111,
    22'b1111111110100011110110,
    22'b1111111111000010100100,
    22'b1111111111100001010010,
    22'b1111111111110101110001,
    22'b0000000000000000000000,
    22'b0000000000001010001111,
    22'b0000000000001010001111,
    22'b0000000000000000000000,
    22'b1111111111110101110001,
    22'b1111111111101011100001,
    22'b1111111111010111000011,
    22'b1111111111000010100100,
    22'b1111111110101110000101,
    22'b1111111110100011110110,
    22'b1111111110001111010111,
    22'b1111111110000101001000,
    22'b1111111110000101001000,
    22'b1111111101111010111000,
    22'b1111111110000101001000,
    22'b1111111110000101001000,
    22'b1111111110001111010111,
    22'b1111111110011001100110,
    22'b1111111110101110000101,
    22'b1111111110111000010100,
    22'b1111111111000010100100,
    22'b1111111111010111000011,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111010111000011,
    22'b1111111111001100110011,
    22'b1111111111001100110011,
    22'b1111111110111000010100,
    22'b1111111110111000010100,
    22'b1111111110111000010100,
    22'b1111111111000010100100,
    22'b1111111111100001010010,
    22'b1111111111010111000011,
    22'b1111111111001100110011,
    22'b0000000000011110101110,
    22'b0000000001010001111011,
    22'b0000000010000101001000,
    22'b0000000011101011100001,
    22'b0000000100011110101110,
    22'b0000000011101011100001,
    22'b0000000001011100001010,
    22'b1111111110001111010111,
    22'b1111111011110101110001,
    22'b1111111010101110000101,
    22'b1111111010101110000101,
    22'b1111111010111000010100,
    22'b1111111010111000010100,
    22'b1111111010000101001000,
    22'b1111111001100110011010,
    22'b1111111001100110011010,
    22'b1111111010011001100110,
    22'b1111111100010100011111,
    22'b1111111101100110011010,
    22'b1111111110101110000101,
    22'b1111111111010111000011,
    22'b1111111111101011100001,
    22'b0000000000000000000000,
    22'b0000000000011110101110,
    22'b0000000000111101011100,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001000111101100,
    22'b0000000000011110101110,
    22'b1111111111100001010010,
    22'b1111111110111000010100,
    22'b1111111110011001100110,
    22'b1111111110000101001000,
    22'b1111111101110000101001,
    22'b1111111100101000111101,
    22'b1111111110100011110110,
    22'b1111111110100011110110,
    22'b1111111011100001010010,
    22'b1111110101110000101001,
    22'b1111110011000010100100,
    22'b1111101101011100001010,
    22'b1111110010011001100110,
    22'b1111110001111010111000,
    22'b1111101110100011110110,
    22'b1111101010011001100110,
    22'b1111100110001111010111,
    22'b1111100011100001010010,
    22'b1111100100111101011100,
    22'b1111100111010111000011,
    22'b1111101011000010100100,
    22'b1111110001010001111011,
    22'b1111111110100011110110,
    22'b0000001000010100011111,
    22'b1111110101111010111000,
    22'b1111110101010001111011,
    22'b1111111001110000101001,
    22'b0000000100101000111101,
    22'b0000010001010001111011,
    22'b0000100011100001010010,
    22'b0000110000001010001111,
    22'b0000110010001111010111,
    22'b0000100011101011100001,
    22'b0000011110111000010100,
    22'b0000010100111101011100,
    22'b0000001011001100110011,
    22'b0000000101010001111011,
    22'b0000000110001111010111,
    22'b1111111110100011110110,
    22'b1111110011010111000011,
    22'b1111100110011001100110,
    22'b1111011100011110101110,
    22'b1111010101110000101001,
    22'b1111010101111010111000,
    22'b1111011010001111010111,
    22'b1111011101011100001010,
    22'b1111100010001111010111,
    22'b1111101000011110101110,
    22'b1111101110000101001000,
    22'b1111110101010001111011,
    22'b1111111110000101001000,
    22'b0000001010100011110110,
    22'b0000010011101011100001,
    22'b0000011011110101110001,
    22'b0000100001111010111000,
    22'b0000100101111010111000,
    22'b0000100010101110000101,
    22'b0000100101000111101100,
    22'b0000100000010100011111,
    22'b0000011001011100001010,
    22'b0000010001000111101100,
    22'b0000001110100011110110,
    22'b0000000111001100110011,
    22'b1111111111110101110001,
    22'b1111111000000000000000,
    22'b1111110010001111010111,
    22'b1111101100111101011100,
    22'b1111101010000101001000,
    22'b1111101000000000000000,
    22'b1111100111001100110011,
    22'b1111100111101011100001,
    22'b1111101000110011001101,
    22'b1111101011100001010010,
    22'b1111101111100001010010,
    22'b1111110100011110101110,
    22'b1111111001110000101001,
    22'b0000000000011110101110,
    22'b0000000101000111101100,
    22'b0000001000111101011100,
    22'b0000001100001010001111,
    22'b0000001110101110000101,
    22'b0000001111000010100100,
    22'b0000001111101011100001,
    22'b0000001101010001111011,
    22'b0000001010000101001000,
    22'b0000001000010100011111,
    22'b0000000101100110011010,
    22'b0000000010100011110110,
    22'b0000000000001010001111,
    22'b1111111100011110101110,
    22'b1111111001100110011010,
    22'b1111110111101011100001,
    22'b1111110110100011110110,
    22'b1111110101100110011010,
    22'b1111110101110000101001,
    22'b1111110110100011110110,
    22'b1111110111010111000011,
    22'b1111111001011100001010,
    22'b1111111011010111000011,
    22'b1111111101011100001010,
    22'b0000000000011110101110,
    22'b0000000010100011110110,
    22'b0000000100011110101110,
    22'b0000000101100110011010,
    22'b0000000110000101001000,
    22'b0000000110011001100110,
    22'b0000000101100110011010,
    22'b0000000100101000111101,
    22'b0000000100000000000000,
    22'b0000000010101110000101,
    22'b0000000001100110011010,
    22'b0000000000001010001111,
    22'b1111111110101110000101,
    22'b1111111101110000101001,
    22'b1111111100101000111101,
    22'b1111111000010100011111,
    22'b1111100000001010001111,
    22'b1111000100010100011111,
    22'b1111100100101000111101,
    22'b1111101101100110011010,
    22'b1111110010100011110110,
    22'b1111110010000101001000,
    22'b1111110110001111010111,
    22'b1111111100111101011100,
    22'b0000010000001010001111,
    22'b0000100000101000111101,
    22'b0000101001100110011010,
    22'b0000101001111010111000,
    22'b0000100110111000010100,
    22'b0000011100110011001101,
    22'b0000011101010001111011,
    22'b0000100101010001111011,
    22'b0000101010001111010111,
    22'b0000101001010001111011,
    22'b0000100101100110011010,
    22'b0000011110011001100110,
    22'b0000010111010111000011,
    22'b0000001110000101001000,
    22'b0000000110111000010100,
    22'b1111111110111000010100,
    22'b1111110111001100110011,
    22'b1111110010100011110110,
    22'b1111110001111010111000,
    22'b1111110010101110000101,
    22'b1111110101010001111011,
    22'b1111111001110000101001,
    22'b1111111100111101011100,
    22'b0000000000000000000000,
    22'b0000000010100011110110,
    22'b0000000100110011001101,
    22'b0000000111100001010010,
    22'b0000001000111101011100,
    22'b0000001001110000101001,
    22'b0000001001100110011010,
    22'b0000000110011001100110,
    22'b0000000011010111000011,
    22'b0000000000001010001111,
    22'b1111111101000111101100,
    22'b1111111001110000101001,
    22'b1111110101111010111000,
    22'b1111110011000010100100,
    22'b1111110000010100011111,
    22'b1111101101011100001010,
    22'b1111101010111000010100,
    22'b1111101001010001111011,
    22'b1111101001010001111011,
    22'b1111101001100110011010,
    22'b1111101000011110101110,
    22'b1111100111100001010010,
    22'b1111100110111000010100,
    22'b1111100110101110000101,
    22'b1111100110100011110110,
    22'b1111100101100110011010,
    22'b1111100100111101011100,
    22'b1111100100000000000000,
    22'b1111100001111010111000,
    22'b1111011111001100110011,
    22'b1111011010011001100110,
    22'b1111010110100011110110,
    22'b1111010011000010100100,
    22'b1111010000011110101110,
    22'b1111001101100110011010,
    22'b1111001011101011100001,
    22'b1111001001011100001010,
    22'b1111000111110101110001,
    22'b1111000101111010111000,
    22'b1111000011100001010010,
    22'b1111000010101110000101,
    22'b1111000010111000010100,
    22'b1111000011100001010010,
    22'b1111000100110011001101,
    22'b1111001011010111000011,
    22'b1111010100111101011100,
    22'b1111011101011100001010,
    22'b1111100001100110011010,
    22'b1111100010100011110110,
    22'b1111011111100001010010,
    22'b1111011011100001010010,
    22'b1111011000000000000000,
    22'b1111010101010001111011,
    22'b1111010000001010001111,
    22'b1111001000010100011111,
    22'b1111000010100011110110,
    22'b1110111001110000101001,
    22'b1110110001111010111000,
    22'b1110101111000010100100,
    22'b1110101100000000000000,
    22'b1110101010011001100110,
    22'b1110101010111000010100,
    22'b1110100111100001010010,
    22'b1110100101110000101001,
    22'b1110100110111000010100,
    22'b1110100111100001010010,
    22'b1110101001000111101100,
    22'b1110101001100110011010,
    22'b1110101101010001111011,
    22'b1110110010111000010100,
    22'b1110110110101110000101,
    22'b1110111011000010100100,
    22'b1110111100001010001111,
    22'b1110110110001111010111,
    22'b1110110011010111000011,
    22'b1110101111100001010010,
    22'b1110101001111010111000,
    22'b1110011100111101011100,
    22'b1110010010111000010100,
    22'b1110010000111101011100,
    22'b1110010001110000101001,
    22'b1110010111101011100001,
    22'b1110111010101110000101,
    22'b1111101000001010001111,
    22'b1111100011101011100001,
    22'b1111011011010111000011,
    22'b1111001100111101011100,
    22'b1110111011101011100001,
    22'b1110111001010001111011,
    22'b1111001101010001111011,
    22'b1111011101100110011010,
    22'b1111100111100001010010,
    22'b1111101010001111010111,
    22'b1111100111001100110011,
    22'b1111011100001010001111,
    22'b1111010001110000101001,
    22'b1111001000111101011100,
    22'b1111000000111101011100,
    22'b1110111000111101011100,
    22'b1110111000001010001111,
    22'b1110111100101000111101,
    22'b1111000100101000111101,
    22'b1111001110000101001000,
    22'b1111011011110101110001,
    22'b1111100110101110000101,
    22'b1111110000000000000000,
    22'b1111110110001111010111,
    22'b1111111000110011001101,
    22'b1111110111000010100100,
    22'b1111110011100001010010,
    22'b1111101111100001010010,
    22'b1111100111110101110001,
    22'b1111011101111010111000,
    22'b1111011000111101011100,
    22'b1111010101111010111000,
    22'b1111010011101011100001,
    22'b1111010000111101011100,
    22'b1111001111101011100001,
    22'b1111010000101000111101,
    22'b1111010011000010100100,
    22'b1111010110000101001000,
    22'b1111011001110000101001,
    22'b1111011011101011100001,
    22'b1111011101100110011010,
    22'b1111011110111000010100,
    22'b1111011111110101110001,
    22'b1111100000000000000000,
    22'b1111011111101011100001,
    22'b1111011111001100110011,
    22'b1111011110111000010100,
    22'b1111011110100011110110,
    22'b1111011101111010111000,
    22'b1111011100111101011100,
    22'b1111011011100001010010,
    22'b1111011001110000101001,
    22'b1111011000110011001101,
    22'b1111011001000111101100,
    22'b1111011001111010111000,
    22'b1111011100000000000000,
    22'b1111011110011001100110,
    22'b1111100001010001111011,
    22'b1111100011100001010010,
    22'b1111100111101011100001,
    22'b1111101010100011110110,
    22'b1111101101100110011010,
    22'b1111110000101000111101,
    22'b1111110101000111101100,
    22'b1111111000010100011111,
    22'b1111111011110101110001,
    22'b1111111111110101110001,
    22'b0000000101100110011010,
    22'b0000001001110000101001,
    22'b0000001100110011001101,
    22'b0000001110001111010111,
    22'b0000001101100110011010,
    22'b0000001010000101001000,
    22'b0000000110000101001000,
    22'b0000000001110000101001,
    22'b1111111101111010111000,
    22'b1111111010000101001000,
    22'b1111111000101000111101,
    22'b1111111000001010001111,
    22'b1111111000011110101110,
    22'b1111111001010001111011,
    22'b1111111010101110000101,
    22'b1111111100000000000000,
    22'b1111111101010001111011,
    22'b1111111110001111010111,
    22'b1111111110111000010100,
    22'b1111111110100011110110,
    22'b1111111101100110011010,
    22'b1111111100101000111101,
    22'b1111111011001100110011,
    22'b1111111010001111010111,
    22'b1111111001010001111011,
    22'b1111111000000000000000,
    22'b1111110110011001100110,
    22'b1111110101000111101100,
    22'b1111110010001111010111,
    22'b1111101010111000010100,
    22'b1111100011110101110001,
    22'b1111011011100001010010,
    22'b1111010001110000101001,
    22'b1111000111010111000011,
    22'b1111000000000000000000,
    22'b1111010100000000000000,
    22'b1111011101010001111011,
    22'b1111100110011001100110,
    22'b1111101010001111010111,
    22'b1111101100101000111101,
    22'b1111101100011110101110,
    22'b1111101010101110000101,
    22'b1111101000110011001101,
    22'b1111100100001010001111,
    22'b1111011000000000000000,
    22'b1111010001100110011010,
    22'b1111001110000101001000,
    22'b1111001100101000111101,
    22'b1111001100110011001101,
    22'b1111001101110000101001,
    22'b1111001111100001010010,
    22'b1111010010001111010111,
    22'b1111010100011110101110,
    22'b1111010101011100001010,
    22'b1111010101111010111000,
    22'b1111010110011001100110,
    22'b1111010110100011110110,
    22'b1111010111000010100100,
    22'b1111010111101011100001,
    22'b1111011000011110101110,
    22'b1111011000011110101110,
    22'b1111011000001010001111,
    22'b1111010111110101110001,
    22'b1111010110101110000101,
    22'b1111010101110000101001,
    22'b1111010100110011001101,
    22'b1111010100000000000000,
    22'b1111010010111000010100,
    22'b1111010001111010111000,
    22'b1111010000110011001101,
    22'b1111010000101000111101,
    22'b1111010001110000101001,
    22'b1111010100111101011100,
    22'b1111011000010100011111,
    22'b1111011100010100011111,
    22'b1111011111110101110001,
    22'b1111100100010100011111,
    22'b1111100111010111000011,
    22'b1111101010100011110110,
    22'b1111101111100001010010,
    22'b1111110011100001010010,
    22'b1111111100110011001101,
    22'b0000000010101110000101,
    22'b0000000111000010100100,
    22'b0000001100011110101110,
    22'b0000010010001111010111,
    22'b0000010010100011110110,
    22'b0000010010111000010100,
    22'b0000010101011100001010,
    22'b0000011001011100001010,
    22'b0000100000110011001101,
    22'b0000100100000000000000,
    22'b0000100011100001010010,
    22'b0000011111100001010010,
    22'b0000010111110101110001,
    22'b0000001011101011100001,
    22'b0000000010101110000101,
    22'b1111111100001010001111,
    22'b1111111000101000111101,
    22'b1111111000111101011100,
    22'b1111111010101110000101,
    22'b1111111100101000111101,
    22'b1111111110001111010111,
    22'b1111111111001100110011,
    22'b1111111111001100110011,
    22'b1111111110101110000101,
    22'b1111111110001111010111,
    22'b1111111110101110000101,
    22'b0000000000111101011100,
    22'b0000000011010111000011,
    22'b0000000101111010111000,
    22'b0000001000010100011111,
    22'b0000001011000010100100,
    22'b0000001100101000111101,
    22'b0000001110100011110110,
    22'b0000010000101000111101,
    22'b0000010001111010111000,
    22'b0000010110001111010111,
    22'b0000011001111010111000,
    22'b0000011001100110011010,
    22'b0000011000011110101110,
    22'b0000011010111000010100,
    22'b0000011000110011001101,
    22'b0000011000010100011111,
    22'b0000011010001111010111,
    22'b0000011001000111101100,
    22'b0000011000001010001111,
    22'b0000010110101110000101,
    22'b0000010100011110101110,
    22'b0000010001110000101001,
    22'b0000001110101110000101,
    22'b0000001100101000111101,
    22'b0000001011010111000011,
    22'b0000001010011001100110,
    22'b0000001001111010111000,
    22'b0000001001011100001010,
    22'b0000001000111101011100,
    22'b0000001000101000111101,
    22'b0000001000011110101110,
    22'b0000000111101011100001,
    22'b0000000111101011100001,
    22'b0000001000010100011111,
    22'b0000001000101000111101,
    22'b0000001001100110011010,
    22'b0000001010100011110110,
    22'b0000001011010111000011,
    22'b0000001100101000111101,
    22'b0000001101000111101100,
    22'b0000001101100110011010,
    22'b0000001101011100001010,
    22'b0000001100011110101110,
    22'b0000001011101011100001,
    22'b0000001010100011110110,
    22'b0000001001010001111011,
    22'b0000001000011110101110,
    22'b0000000111101011100001,
    22'b0000000110111000010100,
    22'b0000000110101110000101,
    22'b0000000110001111010111,
    22'b0000000110011001100110,
    22'b0000000110011001100110,
    22'b0000000101111010111000,
    22'b0000000101100110011010,
    22'b0000000101000111101100,
    22'b0000000100110011001101,
    22'b0000000100110011001101,
    22'b0000000100010100011111,
    22'b0000000100000000000000,
    22'b0000000011101011100001,
    22'b0000000011001100110011,
    22'b0000000010011001100110,
    22'b0000000001100110011010,
    22'b0000000000101000111101,
    22'b1111111111001100110011,
    22'b1111111101010001111011,
    22'b1111111011110101110001,
    22'b1111111010011001100110,
    22'b1111111001010001111011,
    22'b1111111000001010001111,
    22'b1111111000011110101110,
    22'b1111111001111010111000,
    22'b1111111010101110000101,
    22'b1111111100101000111101,
    22'b0000000010100011110110,
    22'b0000000011110101110001,
    22'b0000000010111000010100,
    22'b0000000011001100110011,
    22'b0000000101000111101100,
    22'b0000000101100110011010,
    22'b0000000011110101110001,
    22'b0000000110000101001000,
    22'b0000000110001111010111,
    22'b0000000110100011110110,
    22'b0000001010000101001000,
    22'b0000000101011100001010,
    22'b0000000010101110000101,
    22'b0000000001000111101100,
    22'b1111111111101011100001,
    22'b0000000100000000000000,
    22'b0000001000101000111101,
    22'b0000001000110011001101,
    22'b0000001101110000101001,
    22'b0000010111100001010010,
    22'b0000100000001010001111,
    22'b0000100100101000111101,
    22'b0000101011110101110001,
    22'b0000110010101110000101,
    22'b0000110001111010111000,
    22'b0000101111000010100100,
    22'b0000101011010111000011,
    22'b0000100011001100110011,
    22'b0000010111010111000011,
    22'b0000010010101110000101,
    22'b0000010001110000101001,
    22'b0000010001011100001010,
    22'b0000001010100011110110,
    22'b0000001000011110101110,
    22'b0000001111010111000011,
    22'b0000010100111101011100,
    22'b0000010010001111010111,
    22'b0000011100010100011111,
    22'b1111100100110011001101,
    22'b1110111100011110101110,
    22'b1110111001011100001010,
    22'b1110111000011110101110,
    22'b1110111111000010100100,
    22'b1111000111100001010010,
    22'b1111011001111010111000,
    22'b1111101110111000010100,
    22'b0000001000001010001111,
    22'b0000010010000101001000,
    22'b0000010100101000111101,
    22'b0000010001110000101001,
    22'b0000001101011100001010,
    22'b0000001101010001111011,
    22'b0000001110100011110110,
    22'b0000001101100110011010,
    22'b0000001010011001100110,
    22'b1111011111100001010010,
    22'b1111011110100011110110,
    22'b1111100001010001111011,
    22'b1111101001110000101001,
    22'b1111101111100001010010,
    22'b1111101011010111000011,
    22'b1111011100110011001101,
    22'b1111001001110000101001,
    22'b1111000000010100011111,
    22'b1110110110101110000101,
    22'b1110101101011100001010,
    22'b1110100110000101001000,
    22'b1110101000110011001101,
    22'b1110101011110101110001,
    22'b1110101000010100011111,
    22'b1110011101111010111000,
    22'b1110010110000101001000,
    22'b1110001110000101001000,
    22'b1110000101100110011010,
    22'b1101110100101000111101,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101111000010100011111,
    22'b1110010010111000010100,
    22'b1110100001011100001010,
    22'b1110101001010001111011,
    22'b1110101100110011001101,
    22'b1110101100101000111101,
    22'b1110101010101110000101,
    22'b1110100110011001100110,
    22'b1110100001111010111000,
    22'b1110011011000010100100,
    22'b1110010101110000101001,
    22'b1110001110100011110110,
    22'b1110001010011001100110,
    22'b1110001000010100011111,
    22'b1110001011001100110011,
    22'b1110001011110101110001,
    22'b1110010000001010001111,
    22'b1110010010011001100110,
    22'b1110010110011001100110,
    22'b1110011001100110011010,
    22'b1110011110100011110110,
    22'b1110100101100110011010,
    22'b1110100101100110011010,
    22'b1110100011100001010010,
    22'b1110100010011001100110,
    22'b1110100011110101110001,
    22'b1110100110001111010111,
    22'b1110101000010100011111,
    22'b1110101011010111000011,
    22'b1110101101110000101001,
    22'b1110110011110101110001,
    22'b1110111010011001100110,
    22'b1110111110001111010111,
    22'b1111000100001010001111,
    22'b1111010110001111010111,
    22'b1111011000110011001101,
    22'b1111011001000111101100,
    22'b1111011000111101011100,
    22'b1111011000000000000000,
    22'b1111010110101110000101,
    22'b1111010100011110101110,
    22'b1111010010100011110110,
    22'b1111010000010100011111,
    22'b1111001101011100001010,
    22'b1111001001000111101100,
    22'b1111000101111010111000,
    22'b1111000011001100110011,
    22'b1111000001010001111011,
    22'b1111000000000000000000,
    22'b1110111111010111000011,
    22'b1110111111000010100100,
    22'b1110111111000010100100,
    22'b1110111110111000010100,
    22'b1110111110111000010100,
    22'b1110111111010111000011,
    22'b1110111111110101110001,
    22'b1110111110101110000101,
    22'b1111000001000111101100,
    22'b1111000011010111000011,
    22'b1111000100011110101110,
    22'b1111000101100110011010,
    22'b1111000110111000010100,
    22'b1111001000010100011111,
    22'b1111001010111000010100,
    22'b1111001101011100001010,
    22'b1111001101110000101001,
    22'b1111001101111010111000,
    22'b1111001111100001010010,
    22'b1111010001000111101100,
    22'b1111010010111000010100,
    22'b1111010100110011001101,
    22'b1111010111000010100100,
    22'b1111011000111101011100,
    22'b1111011011100001010010,
    22'b1111011101110000101001,
    22'b1111100101011100001010,
    22'b1111101100011110101110,
    22'b1111110001100110011010,
    22'b1111111000000000000000,
    22'b0000000000000000000000,
    22'b0000000011101011100001,
    22'b0000000110101110000101,
    22'b0000001110111000010100,
    22'b0000010001011100001010,
    22'b0000010100010100011111,
    22'b0000010111010111000011,
    22'b0000011001011100001010,
    22'b0000011001111010111000,
    22'b0000011100010100011111,
    22'b0000011110111000010100,
    22'b0000011101100110011010,
    22'b0000011111010111000011,
    22'b0000011111110101110001,
    22'b0000100001000111101100,
    22'b0000100010001111010111,
    22'b0000100100011110101110,
    22'b0000100101000111101100,
    22'b0000100101111010111000,
    22'b0000100111000010100100,
    22'b0000101000101000111101,
    22'b0000101001111010111000,
    22'b0000101011101011100001,
    22'b0000101101011100001010,
    22'b0000101110111000010100,
    22'b0000110000110011001101,
    22'b0000110010011001100110,
    22'b0000110010101110000101,
    22'b0000110100111101011100,
    22'b0000111001010001111011,
    22'b0000111110100011110110,
    22'b0001000100111101011100,
    22'b0001001000010100011111,
    22'b0001001010100011110110,
    22'b0001001011000010100100,
    22'b0001001010011001100110,
    22'b0001001011001100110011,
    22'b0001001101100110011010,
    22'b0001010000110011001101,
    22'b0001010100010100011111,
    22'b0001011000000000000000,
    22'b0001011100011110101110,
    22'b0001011110111000010100,
    22'b0001100000000000000000,
    22'b0001100000111101011100,
    22'b0001100010100011110110,
    22'b0001100100010100011111,
    22'b0001100110100011110110,
    22'b0001101001011100001010,
    22'b0001101101000111101100,
    22'b0001110011010111000011,
    22'b0001111000000000000000,
    22'b0001111011100001010010,
    22'b0010000010000101001000,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011010111000011,
    22'b0010001011100001010010,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001011101011100001,
    22'b0010001000110011001101,
    22'b0010000100011110101110,
    22'b0001111100011110101110,
    22'b0001110100001010001111,
    22'b0001101010001111010111,
    22'b0001100000110011001101,
    22'b0001010111010111000011,
    22'b0001010001111010111000,
    22'b0001001110000101001000,
    22'b0001001110011001100110,
    22'b0001001100010100011111,
    22'b0001001010001111010111,
    22'b0001000110000101001000,
    22'b0001000000101000111101,
    22'b0000111011000010100100,
    22'b0000110110100011110110,
    22'b0000110101000111101100,
    22'b0000110100000000000000,
    22'b0000110010111000010100,
    22'b0000110001010001111011,
    22'b0000110000000000000000,
    22'b0000101110101110000101,
    22'b0000101110000101001000,
    22'b0000101101111010111000,
    22'b0000101101100110011010,
    22'b0000101100101000111101,
    22'b0000101011110101110001,
    22'b0000101011010111000011,
    22'b0000101010111000010100,
    22'b0000101001110000101001,
    22'b0000101000011110101110,
    22'b0000100110101110000101,
    22'b0000100100101000111101,
    22'b0000100100110011001101,
    22'b0000100111001100110011,
    22'b0000101001100110011010,
    22'b0000101010000101001000,
    22'b0000100111110101110001,
    22'b0000100100011110101110,
    22'b0000100001110000101001,
    22'b0000100000001010001111,
    22'b0000100000111101011100,
    22'b0000011111010111000011,
    22'b0000011101111010111000,
    22'b0000011100000000000000,
    22'b0000011011100001010010,
    22'b0000011010001111010111,
    22'b0000011000011110101110,
    22'b0000010101011100001010,
    22'b0000010011100001010010,
    22'b0000010000111101011100,
    22'b0000001100011110101110,
    22'b0000000011010111000011,
    22'b1111111010011001100110,
    22'b1111110000101000111101,
    22'b1111100111100001010010,
    22'b1111010011101011100001,
    22'b1111010010100011110110,
    22'b1111010000111101011100,
    22'b1111001101100110011010,
    22'b1111000111100001010010,
    22'b1110111011101011100001,
    22'b1110101100000000000000,
    22'b1110011110011001100110,
    22'b1110001110100011110110,
    22'b1110000100101000111101,
    22'b1101111101010001111011,
    22'b1101111011110101110001,
    22'b1101111110001111010111,
    22'b1110000010011001100110,
    22'b1110000110101110000101,
    22'b1110001001010001111011,
    22'b1110001010000101001000,
    22'b1110001100110011001101,
    22'b1110010110011001100110,
    22'b1110100010011001100110,
    22'b1110101111110101110001,
    22'b1111000001111010111000,
    22'b1111001101011100001010,
    22'b1111010101100110011010,
    22'b1111011010000101001000,
    22'b1111011011001100110011,
    22'b1111011010001111010111,
    22'b1111011001011100001010,
    22'b1111011001000111101100,
    22'b1111011101110000101001,
    22'b1111100010001111010111,
    22'b1111011111001100110011,
    22'b1111010100101000111101,
    22'b1111000101000111101100,
    22'b1110111011100001010010,
    22'b1110110100110011001101,
    22'b1110110010000101001000,
    22'b1110100100111101011100,
    22'b1110000011000010100100,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110100010100011111,
    22'b1101110110100011110110,
    22'b1101111000000000000000,
    22'b1101111000110011001101,
    22'b1101111011000010100100,
    22'b1101111100011110101110,
    22'b1101111101011100001010,
    22'b1101111101110000101001,
    22'b1101111101100110011010,
    22'b1101111101010001111011,
    22'b1101111101110000101001,
    22'b1101111111110101110001,
    22'b1110000110001111010111,
    22'b1110001011110101110001,
    22'b1110010000010100011111,
    22'b1110010011001100110011,
    22'b1110010100101000111101,
    22'b1110010100101000111101,
    22'b1110010100010100011111,
    22'b1110010100011110101110,
    22'b1110010101100110011010,
    22'b1110011000011110101110,
    22'b1110011011010111000011,
    22'b1110011110101110000101,
    22'b1110100001111010111000,
    22'b1110100101110000101001,
    22'b1110101000001010001111,
    22'b1110101010001111010111,
    22'b1110101011110101110001,
    22'b1110101101111010111000,
    22'b1110101110111000010100,
    22'b1110101111001100110011,
    22'b1110101110101110000101,
    22'b1110101101010001111011,
    22'b1110101011000010100100,
    22'b1110101001011100001010,
    22'b1110101000011110101110,
    22'b1110101000011110101110,
    22'b1110101001100110011010,
    22'b1110101011000010100100,
    22'b1110101100010100011111,
    22'b1110101100110011001101,
    22'b1110101100010100011111,
    22'b1110101011101011100001,
    22'b1110101011000010100100,
    22'b1110101011000010100100,
    22'b1110101011110101110001,
    22'b1110101110000101001000,
    22'b1110110000001010001111,
    22'b1110110010000101001000,
    22'b1110110011101011100001,
    22'b1110110101011100001010,
    22'b1110110110001111010111,
    22'b1110110101010001111011,
    22'b1110110111001100110011,
    22'b1110111010011001100110,
    22'b1110111100010100011111,
    22'b1110111101011100001010,
    22'b1110111111100001010010,
    22'b1110111111100001010010,
    22'b1110111110111000010100,
    22'b1110111101000111101100,
    22'b1110111000010100011111,
    22'b1110110011101011100001,
    22'b1110101110100011110110,
    22'b1110101001100110011010,
    22'b1110100100001010001111,
    22'b1110100001010001111011,
    22'b1110011111101011100001,
    22'b1110011111100001010010,
    22'b1110100000110011001101,
    22'b1110100010100011110110,
    22'b1110100100011110101110,
    22'b1110100101110000101001,
    22'b1110100110001111010111,
    22'b1110100110011001100110,
    22'b1110100110101110000101,
    22'b1110100111100001010010,
    22'b1110101001011100001010,
    22'b1110101011100001010010,
    22'b1110101110000101001000,
    22'b1110110010011001100110,
    22'b1110111011010111000011,
    22'b1111000010011001100110,
    22'b1111000111010111000011,
    22'b1111001001100110011010,
    22'b1111001010011001100110,
    22'b1111001011000010100100,
    22'b1111001100001010001111,
    22'b1111001101111010111000,
    22'b1111010000101000111101,
    22'b1111010100111101011100,
    22'b1111011000011110101110,
    22'b1111011100010100011111,
    22'b1111100000111101011100,
    22'b1111100100001010001111,
    22'b1111100111100001010010,
    22'b1111101011000010100100,
    22'b1111101111101011100001,
    22'b1111110010101110000101,
    22'b1111110101011100001010,
    22'b1111111000000000000000,
    22'b1111111011000010100100,
    22'b0000000000001010001111,
    22'b0000000100011110101110,
    22'b0000001001000111101100,
    22'b0000001101110000101001,
    22'b0000010011101011100001,
    22'b0000011000001010001111,
    22'b0000011100001010001111,
    22'b0000011111101011100001,
    22'b0000100011110101110001,
    22'b0000100110100011110110,
    22'b0000101000110011001101,
    22'b0000101010101110000101,
    22'b0000101100101000111101,
    22'b0000101111010111000011,
    22'b0000110001111010111000,
    22'b0000110100101000111101,
    22'b0000110111110101110001,
    22'b0000111011110101110001,
    22'b0000111110011001100110,
    22'b0001000000101000111101,
    22'b0001000010000101001000,
    22'b0001000010011001100110,
    22'b0001000010001111010111,
    22'b0001000001110000101001,
    22'b0001000001010001111011,
    22'b0001000000110011001101,
    22'b0001000001010001111011,
    22'b0001000010100011110110,
    22'b0001000100001010001111,
    22'b0001000110001111010111,
    22'b0001001010000101001000,
    22'b0001001110000101001000,
    22'b0001010001100110011010,
    22'b0001010100110011001101,
    22'b0001011010000101001000,
    22'b0001101000001010001111,
    22'b0001101111010111000011,
    22'b0001110011100001010010,
    22'b0001110010101110000101,
    22'b0001101101000111101100,
    22'b0001101000101000111101,
    22'b0001100011010111000011,
    22'b0001011101100110011010,
    22'b0001010111001100110011,
    22'b0001001001111010111000,
    22'b0001000010101110000101,
    22'b0000111110101110000101,
    22'b0000111100010100011111,
    22'b0000111011000010100100,
    22'b0000111011010111000011,
    22'b0000111100000000000000,
    22'b0000111101000111101100,
    22'b0000111110001111010111,
    22'b0000111111010111000011,
    22'b0001000000011110101110,
    22'b0001000001100110011010,
    22'b0001000010111000010100,
    22'b0001000100110011001101,
    22'b0001001010000101001000,
    22'b0001010010000101001000,
    22'b0001011010000101001000,
    22'b0001011111001100110011,
    22'b0001100100010100011111,
    22'b0001100100000000000000,
    22'b0001100000111101011100,
    22'b0001011101111010111000,
    22'b0001011010101110000101,
    22'b0001011000101000111101,
    22'b0001010110101110000101,
    22'b0001010010100011110110,
    22'b0001001100111101011100,
    22'b0001000110000101001000,
    22'b0000111110100011110110,
    22'b0000111100111101011100,
    22'b0000111100101000111101,
    22'b0000111011101011100001,
    22'b0000111010100011110110,
    22'b0000111001110000101001,
    22'b0000111000000000000000,
    22'b0000110101100110011010,
    22'b0000110011001100110011,
    22'b0000110000011110101110,
    22'b0000101100111101011100,
    22'b0000101010111000010100,
    22'b0000101000111101011100,
    22'b0000100111100001010010,
    22'b0000100110111000010100,
    22'b0000100111001100110011,
    22'b0000100111110101110001,
    22'b0000101010000101001000,
    22'b0000101101111010111000,
    22'b0000110010111000010100,
    22'b0000110101111010111000,
    22'b0000111010001111010111,
    22'b0000111110011001100110,
    22'b0001000100010100011111,
    22'b0001001000111101011100,
    22'b0001001001011100001010,
    22'b0001000100011110101110,
    22'b0000111101011100001010,
    22'b0000110110101110000101,
    22'b0000110010101110000101,
    22'b0000110010000101001000,
    22'b0000110100111101011100,
    22'b0000111010011001100110,
    22'b0001000011101011100001,
    22'b0001001000001010001111,
    22'b0001001001100110011010,
    22'b0001000100010100011111,
    22'b0000111100010100011111,
    22'b0000101110000101001000,
    22'b0000100011001100110011,
    22'b0000011001111010111000,
    22'b0000010011000010100100,
    22'b0000001110011001100110,
    22'b0000001011100001010010,
    22'b0000001011010111000011,
    22'b0000001100001010001111,
    22'b0000001101110000101001,
    22'b0000001111101011100001,
    22'b0000010010011001100110,
    22'b0000010100011110101110,
    22'b0000010110011001100110,
    22'b0000011000010100011111,
    22'b0000011010001111010111,
    22'b0000011101000111101100,
    22'b0000011111001100110011,
    22'b0000100001010001111011,
    22'b0000100011010111000011,
    22'b0000100101010001111011,
    22'b0000100111100001010010,
    22'b0000101000101000111101,
    22'b0000101001010001111011,
    22'b0000101001011100001010,
    22'b0000101001000111101100,
    22'b0000100111110101110001,
    22'b0000100110011001100110,
    22'b0000100100101000111101,
    22'b0000100010101110000101,
    22'b0000100000011110101110,
    22'b0000011111001100110011,
    22'b0000011110100011110110,
    22'b0000011110000101001000,
    22'b0000011110001111010111,
    22'b0000011110101110000101,
    22'b0000011111100001010010,
    22'b0000100000110011001101,
    22'b0000100010100011110110,
    22'b0000100101110000101001,
    22'b0000101000101000111101,
    22'b0000101100000000000000,
    22'b0000101111001100110011,
    22'b0000110010001111010111,
    22'b0000110101100110011010,
    22'b0000110111010111000011,
    22'b0000110111110101110001,
    22'b0000111000001010001111,
    22'b0000111000000000000000,
    22'b0000111000000000000000,
    22'b0000110111110101110001,
    22'b0000110110101110000101,
    22'b0000110100001010001111,
    22'b0000110000110011001101,
    22'b0000101110011001100110,
    22'b0000101011101011100001,
    22'b0000101001111010111000,
    22'b0000101000010100011111,
    22'b0000100110011001100110,
    22'b0000100100101000111101,
    22'b0000100011010111000011,
    22'b0000100001111010111000,
    22'b0000100000011110101110,
    22'b0000011111000010100100,
    22'b0000011101011100001010,
    22'b0000011100011110101110,
    22'b0000011011101011100001,
    22'b0000011011000010100100,
    22'b0000011011000010100100,
    22'b0000011011101011100001,
    22'b0000011100110011001101,
    22'b0000011101111010111000,
    22'b0000011111010111000011,
    22'b0000100001000111101100,
    22'b0000100001110000101001,
    22'b0000100001100110011010,
    22'b0000100000001010001111,
    22'b0000011110000101001000,
    22'b0000011010100011110110,
    22'b0000010111010111000011,
    22'b0000010100011110101110,
    22'b0000010010011001100110,
    22'b0000010000111101011100,
    22'b0000001111001100110011,
    22'b0000001110000101001000,
    22'b0000001100111101011100,
    22'b0000001100000000000000,
    22'b0000001010111000010100,
    22'b0000001001000111101100,
    22'b0000000111100001010010,
    22'b0000000110001111010111,
    22'b0000000101011100001010,
    22'b0000000101011100001010,
    22'b0000000110111000010100,
    22'b0000001001000111101100,
    22'b0000001100001010001111,
    22'b0000001111101011100001,
    22'b0000010011010111000011,
    22'b0000011000010100011111,
    22'b0000011011100001010010,
    22'b0000011110000101001000,
    22'b0000011111100001010010,
    22'b0000011111110101110001,
    22'b0000011111010111000011,
    22'b0000011100111101011100,
    22'b0000011010101110000101,
    22'b0000011000010100011111,
    22'b0000010011110101110001,
    22'b0000010000111101011100,
    22'b0000001101110000101001,
    22'b0000001010001111010111,
    22'b0000000111010111000011,
    22'b0000000100000000000000,
    22'b0000000010000101001000,
    22'b0000000000101000111101,
    22'b1111111111010111000011,
    22'b1111111110100011110110,
    22'b1111111110101110000101,
    22'b0000000000110011001101,
    22'b0000000000111101011100,
    22'b1111111110001111010111,
    22'b1111111010000101001000,
    22'b1111110111010111000011,
    22'b1111110101010001111011,
    22'b1111110011010111000011,
    22'b1111110001100110011010,
    22'b1111110001010001111011,
    22'b1111110001111010111000,
    22'b1111110011000010100100,
    22'b1111110011110101110001,
    22'b1111110100011110101110,
    22'b1111110100010100011111,
    22'b1111110011101011100001,
    22'b1111110010001111010111,
    22'b1111101111101011100001,
    22'b1111101101100110011010,
    22'b1111101011110101110001,
    22'b1111101011100001010010,
    22'b1111101001110000101001,
    22'b1111100110101110000101,
    22'b1111100100011110101110,
    22'b1111100011010111000011,
    22'b1111100010111000010100,
    22'b1111100001100110011010,
    22'b1111011111100001010010,
    22'b1111011100001010001111,
    22'b1111010111101011100001,
    22'b1111010010100011110110,
    22'b1111001011010111000011,
    22'b1111000110100011110110,
    22'b1111000010000101001000,
    22'b1110111111110101110001,
    22'b1110111110101110000101,
    22'b1110111110111000010100,
    22'b1110111111100001010010,
    22'b1111000000000000000000,
    22'b1111000001110000101001,
    22'b1111000100010100011111,
    22'b1111000110100011110110,
    22'b1111001000001010001111,
    22'b1111001000111101011100,
    22'b1111001000101000111101,
    22'b1111001000101000111101,
    22'b1111001000010100011111,
    22'b1111000111100001010010,
    22'b1111000110100011110110,
    22'b1111000110011001100110,
    22'b1111000111000010100100,
    22'b1111001000000000000000,
    22'b1111001000011110101110,
    22'b1111001010011001100110,
    22'b1111001100010100011111,
    22'b1111001111000010100100,
    22'b1111010011010111000011,
    22'b1111010111100001010010,
    22'b1111011011101011100001,
    22'b1111011111101011100001,
    22'b1111100010101110000101,
    22'b1111100100110011001101,
    22'b1111100101000111101100,
    22'b1111100100001010001111,
    22'b1111100010100011110110,
    22'b1111011111101011100001,
    22'b1111011101100110011010,
    22'b1111011011101011100001,
    22'b1111011010011001100110,
    22'b1111011001111010111000,
    22'b1111011010111000010100,
    22'b1111011100111101011100,
    22'b1111100000000000000000,
    22'b1111100011101011100001,
    22'b1111101000111101011100,
    22'b1111101100111101011100,
    22'b1111110000110011001101,
    22'b1111110100011110101110,
    22'b1111111000000000000000,
    22'b1111111100010100011111,
    22'b1111111111001100110011,
    22'b0000000001111010111000,
    22'b0000000100001010001111,
    22'b0000000101111010111000,
    22'b0000001000000000000000,
    22'b0000001001011100001010,
    22'b0000001011101011100001,
    22'b0000001110111000010100,
    22'b0000010000111101011100,
    22'b0000001101111010111000,
    22'b0000000111101011100001,
    22'b0000000000000000000000,
    22'b1111111000010100011111,
    22'b1111110001000111101100,
    22'b1111101010000101001000,
    22'b1111100111101011100001,
    22'b1111101000011110101110,
    22'b1111101100010100011111,
    22'b1111110100011110101110,
    22'b1111111011101011100001,
    22'b0000000010100011110110,
    22'b0000001000111101011100,
    22'b0000001110011001100110,
    22'b0000010100011110101110,
    22'b0000011000101000111101,
    22'b0000011011110101110001,
    22'b0000011110001111010111,
    22'b0000011111101011100001,
    22'b0000100001011100001010,
    22'b0000100010100011110110,
    22'b0000100110101110000101,
    22'b0000101111001100110011,
    22'b0000111010001111010111,
    22'b0001000011101011100001,
    22'b0001000101000111101100,
    22'b0001000010011001100110,
    22'b0000111101000111101100,
    22'b0000110011010111000011,
    22'b0000101101011100001010,
    22'b0000101001100110011010,
    22'b0000100111101011100001,
    22'b0000100111100001010010,
    22'b0000101001100110011010,
    22'b0000101101000111101100,
    22'b0000101101011100001010,
    22'b0000101011010111000011,
    22'b0000100111110101110001,
    22'b0000100010001111010111,
    22'b0000011100001010001111,
    22'b0000010100110011001101,
    22'b0000010000010100011111,
    22'b0000001101000111101100,
    22'b0000001001000111101100,
    22'b0000000101011100001010,
    22'b0000000000111101011100,
    22'b1111111100111101011100,
    22'b1111111000110011001101,
    22'b1111110101111010111000,
    22'b1111110011000010100100,
    22'b1111110000001010001111,
    22'b1111101101011100001010,
    22'b1111101001110000101001,
    22'b1111101000000000000000,
    22'b1111100111001100110011,
    22'b1111100110111000010100,
    22'b1111100111000010100100,
    22'b1111100111001100110011,
    22'b1111100111001100110011,
    22'b1111100111100001010010,
    22'b1111101000001010001111,
    22'b1111100111110101110001,
    22'b1111100110100011110110,
    22'b1111100100111101011100,
    22'b1111100100011110101110,
    22'b1111100101011100001010,
    22'b1111100101100110011010,
    22'b1111100100101000111101,
    22'b1111100100110011001101,
    22'b1111101000011110101110,
    22'b1111101101010001111011,
    22'b1111110010011001100110,
    22'b1111110110101110000101,
    22'b1111111010111000010100,
    22'b1111111100011110101110,
    22'b1111111100111101011100,
    22'b1111111100000000000000,
    22'b1111111000011110101110,
    22'b1111110100011110101110,
    22'b1111101111100001010010,
    22'b1111101010001111010111,
    22'b1111100011001100110011,
    22'b1111011110100011110110,
    22'b1111011010111000010100,
    22'b1111011000011110101110,
    22'b1111010110101110000101,
    22'b1111010101111010111000,
    22'b1111010100110011001101,
    22'b1111011000001010001111,
    22'b1111011011100001010010,
    22'b1111011100101000111101,
    22'b1111011110011001100110,
    22'b1111100100011110101110,
    22'b1111101010100011110110,
    22'b1111101111110101110001,
    22'b1111110010101110000101,
    22'b1111110101000111101100,
    22'b1111110110101110000101,
    22'b1111110101110000101001,
    22'b1111110001111010111000,
    22'b1111101100011110101110,
    22'b1111100101010001111011,
    22'b1111011111110101110001,
    22'b1111011010101110000101,
    22'b1111010110011001100110,
    22'b1111010001100110011010,
    22'b1111001111010111000011,
    22'b1111001100111101011100,
    22'b1111000111010111000011,
    22'b1110111100011110101110,
    22'b1110110011000010100100,
    22'b1110101010000101001000,
    22'b1110100010111000010100,
    22'b1110011110001111010111,
    22'b1110011101010001111011,
    22'b1110011101111010111000,
    22'b1110100000010100011111,
    22'b1110100001000111101100,
    22'b1110100100001010001111,
    22'b1110101000111101011100,
    22'b1110101100000000000000,
    22'b1110101111000010100100,
    22'b1110110010000101001000,
    22'b1110110100110011001101,
    22'b1110110111001100110011,
    22'b1110111010011001100110,
    22'b1110111101000111101100,
    22'b1111000000101000111101,
    22'b1111000100001010001111,
    22'b1111000111101011100001,
    22'b1111001001010001111011,
    22'b1111001010101110000101,
    22'b1111001100010100011111,
    22'b1111001110100011110110,
    22'b1111010000011110101110,
    22'b1111010010100011110110,
    22'b1111010111001100110011,
    22'b1111010110111000010100,
    22'b1111010110000101001000,
    22'b1111010101011100001010,
    22'b1111010100011110101110,
    22'b1111010011101011100001,
    22'b1111010010100011110110,
    22'b1111010001011100001010,
    22'b1111001111100001010010,
    22'b1111001101011100001010,
    22'b1111001010111000010100,
    22'b1111000111110101110001,
    22'b1111000010011001100110,
    22'b1110111101010001111011,
    22'b1110110111100001010010,
    22'b1110101111010111000011,
    22'b1110101001010001111011,
    22'b1110100100011110101110,
    22'b1110100001010001111011,
    22'b1110100000110011001101,
    22'b1110100001111010111000,
    22'b1110100011100001010010,
    22'b1110100101000111101100,
    22'b1110100111010111000011,
    22'b1110101001010001111011,
    22'b1110101011010111000011,
    22'b1110101101000111101100,
    22'b1110101110001111010111,
    22'b1110101110101110000101,
    22'b1110101111101011100001,
    22'b1110110001000111101100,
    22'b1110110011100001010010,
    22'b1110110110001111010111,
    22'b1110111011110101110001,
    22'b1111000010111000010100,
    22'b1111001100000000000000,
    22'b1111010010000101001000,
    22'b1111010110100011110110,
    22'b1111011001010001111011,
    22'b1111011010000101001000,
    22'b1111011001111010111000,
    22'b1111011000011110101110,
    22'b1111010100111101011100,
    22'b1111010001010001111011,
    22'b1111001101011100001010,
    22'b1111001001111010111000,
    22'b1111000101111010111000,
    22'b1111000010101110000101,
    22'b1110111111010111000011,
    22'b1110111011100001010010,
    22'b1110110110011001100110,
    22'b1110110011010111000011,
    22'b1110110001000111101100,
    22'b1110101111100001010010,
    22'b1110101111010111000011,
    22'b1110110000011110101110,
    22'b1110110010001111010111,
    22'b1110110101100110011010,
    22'b1110111000101000111101,
    22'b1110111011110101110001,
    22'b1110111110111000010100,
    22'b1111000001111010111000,
    22'b1111000011101011100001,
    22'b1111000101000111101100,
    22'b1111000110000101001000,
    22'b1111000111001100110011,
    22'b1111000111100001010010,
    22'b1111000111101011100001,
    22'b1111001000010100011111,
    22'b1111001000101000111101,
    22'b1111001000101000111101,
    22'b1111001000011110101110,
    22'b1111000111110101110001,
    22'b1111000111001100110011,
    22'b1111000110111000010100,
    22'b1111000110101110000101,
    22'b1111000111000010100100,
    22'b1111000111110101110001,
    22'b1111001001000111101100,
    22'b1111001011010111000011,
    22'b1111001100111101011100,
    22'b1111001110100011110110,
    22'b1111001111010111000011,
    22'b1111001111001100110011,
    22'b1111001110101110000101,
    22'b1111001110011001100110,
    22'b1111001110011001100110,
    22'b1111001110101110000101,
    22'b1111010000001010001111,
    22'b1111010001100110011010,
    22'b1111010011001100110011,
    22'b1111010100110011001101,
    22'b1111010111001100110011,
    22'b1111011000111101011100,
    22'b1111011011000010100100,
    22'b1111011100111101011100,
    22'b1111011111000010100100,
    22'b1111011111110101110001,
    22'b1111011111110101110001,
    22'b1111011111010111000011,
    22'b1111011110101110000101,
    22'b1111011110001111010111,
    22'b1111011101100110011010,
    22'b1111011100011110101110,
    22'b1111011010111000010100,
    22'b1111011001111010111000,
    22'b1111011001011100001010,
    22'b1111011001011100001010,
    22'b1111011010011001100110,
    22'b1111011011010111000011,
    22'b1111011100010100011111,
    22'b1111011101010001111011,
    22'b1111011110111000010100,
    22'b1111100000000000000000,
    22'b1111100001011100001010,
    22'b1111100011010111000011,
    22'b1111100100110011001101,
    22'b1111100110100011110110,
    22'b1111101000011110101110,
    22'b1111110001000111101100,
    22'b1111110010100011110110,
    22'b1111110100000000000000,
    22'b1111110101011100001010,
    22'b1111110111000010100100,
    22'b1111111000010100011111,
    22'b1111111001110000101001,
    22'b1111111011001100110011,
    22'b1111111100111101011100,
    22'b1111111111100001010010,
    22'b0000000001011100001010,
    22'b0000000011100001010010,
    22'b0000000101100110011010,
    22'b0000001000010100011111,
    22'b0000001010001111010111,
    22'b0000001100001010001111,
    22'b0000001110011001100110,
    22'b0000010000101000111101,
    22'b0000010100000000000000,
    22'b0000010110100011110110,
    22'b0000011001011100001010,
    22'b0000011100000000000000,
    22'b0000011100110011001101,
    22'b0000011010101110000101,
    22'b0000011010101110000101,
    22'b0000011100111101011100,
    22'b0000100000101000111101,
    22'b0000100110000101001000,
    22'b0000101001011100001010,
    22'b0000101100010100011111,
    22'b0000101111000010100100,
    22'b0000110001111010111000,
    22'b0000110011001100110011,
    22'b0000110100010100011111,
    22'b0000110101010001111011,
    22'b0000110110000101001000,
    22'b0000110110101110000101,
    22'b0000110110111000010100,
    22'b0000110111000010100100,
    22'b0000110111001100110011,
    22'b0000111000000000000000,
    22'b0000111000101000111101,
    22'b0000111000010100011111,
    22'b0000110111101011100001,
    22'b0000110110111000010100,
    22'b0000110101011100001010,
    22'b0000110100000000000000,
    22'b0000110011010111000011,
    22'b0000110010101110000101,
    22'b0000110010111000010100,
    22'b0000110101000111101100,
    22'b0000110110111000010100,
    22'b0000111000111101011100,
    22'b0000111011010111000011,
    22'b0001000001111010111000,
    22'b0001000110111000010100,
    22'b0001001011000010100100,
    22'b0001010010101110000101,
    22'b0001100001000111101100,
    22'b0001110110100011110110,
    22'b0001111010000101001000,
    22'b0001110011001100110011,
    22'b0001101010001111010111,
    22'b0001100011001100110011,
    22'b0001011101110000101001,
    22'b0001011011001100110011,
    22'b0001011000001010001111,
    22'b0001010100000000000000,
    22'b0001001111000010100100,
    22'b0001000111001100110011,
    22'b0001000001010001111011,
    22'b0000111011000010100100,
    22'b0000110101110000101001,
    22'b0000101111010111000011,
    22'b0000101011000010100100,
    22'b0000100111000010100100,
    22'b0000100011101011100001,
    22'b0000100000101000111101,
    22'b0000011101011100001010,
    22'b0000011011010111000011,
    22'b0000011001111010111000,
    22'b0000011000110011001101,
    22'b0000011000000000000000,
    22'b0000010101110000101001,
    22'b0000010011110101110001,
    22'b0000011001010001111011,
    22'b0000101001010001111011,
    22'b0000110001100110011010,
    22'b0000101010000101001000,
    22'b0000100000000000000000,
    22'b0000011000110011001101,
    22'b0000010100101000111101,
    22'b0000001110111000010100,
    22'b0000001000110011001101,
    22'b0000000010101110000101,
    22'b1111111110000101001000,
    22'b1111111010000101001000,
    22'b1111110110000101001000,
    22'b1111110001000111101100,
    22'b1111101011001100110011,
    22'b1111011110011001100110,
    22'b1111010010011001100110,
    22'b1111000110111000010100,
    22'b1110111100011110101110,
    22'b1110110001110000101001,
    22'b1110101100011110101110,
    22'b1110101001010001111011,
    22'b1110101000111101011100,
    22'b1110101100001010001111,
    22'b1110101101100110011010,
    22'b1110110001110000101001,
    22'b1110110101011100001010,
    22'b1110110101100110011010,
    22'b1110110011001100110011,
    22'b1110110001100110011010,
    22'b1110110001110000101001,
    22'b1110110011000010100100,
    22'b1110110100011110101110,
    22'b1110110110011001100110,
    22'b1110111000010100011111,
    22'b1110110101000111101100,
    22'b1110110011101011100001,
    22'b1110110001110000101001,
    22'b1110110001100110011010,
    22'b1110101101100110011010,
    22'b1110101100001010001111,
    22'b1110101101110000101001,
    22'b1110110001011100001010,
    22'b1110110110101110000101,
    22'b1110111010011001100110,
    22'b1110111100001010001111,
    22'b1110111101010001111011,
    22'b1110110111000010100100,
    22'b1110110010111000010100,
    22'b1110101110101110000101,
    22'b1110101000110011001101,
    22'b1110100100101000111101,
    22'b1110100000111101011100,
    22'b1110011100011110101110,
    22'b1110011001011100001010,
    22'b1110010110111000010100,
    22'b1110010100110011001101,
    22'b1110010011010111000011,
    22'b1110010011010111000011,
    22'b1110010100010100011111,
    22'b1110010110001111010111,
    22'b1110011001110000101001,
    22'b1110011100110011001101,
    22'b1110100000000000000000,
    22'b1110100011000010100100,
    22'b1110100110101110000101,
    22'b1110101000111101011100,
    22'b1110101010101110000101,
    22'b1110101100011110101110,
    22'b1110101110101110000101,
    22'b1110110000011110101110,
    22'b1110110010001111010111,
    22'b1110110100001010001111,
    22'b1110110111000010100100,
    22'b1110111001000111101100,
    22'b1110111011000010100100,
    22'b1110111100111101011100,
    22'b1110111111110101110001,
    22'b1111000001110000101001,
    22'b1111000011010111000011,
    22'b1111000110001111010111,
    22'b1111001000101000111101,
    22'b1111001010101110000101,
    22'b1111001100110011001101,
    22'b1111001111010111000011,
    22'b1111010000111101011100,
    22'b1111010010100011110110,
    22'b1111010011110101110001,
    22'b1111010101010001111011,
    22'b1111010110011001100110,
    22'b1111010111010111000011,
    22'b1111011000010100011111,
    22'b1111011010001111010111,
    22'b1111011011101011100001,
    22'b1111011100111101011100,
    22'b1111011111001100110011,
    22'b1111100010100011110110,
    22'b1111100100011110101110,
    22'b1111100110011001100110,
    22'b1111101000110011001101,
    22'b1111101100001010001111,
    22'b1111101110001111010111,
    22'b1111101111110101110001,
    22'b1111110001000111101100,
    22'b1111110010011001100110,
    22'b1111110011101011100001,
    22'b1111110101011100001010,
    22'b1111111001011100001010,
    22'b1111111100011110101110,
    22'b1111111111010111000011,
    22'b0000000010001111010111,
    22'b0000010010111000010100,
    22'b0000011000010100011111,
    22'b0000011101111010111000,
    22'b0000101001000111101100,
    22'b0000111001111010111000,
    22'b0001000010001111010111,
    22'b0001001000111101011100,
    22'b0001010000000000000000,
    22'b0001011110001111010111,
    22'b0001100101000111101100,
    22'b0001101010011001100110,
    22'b0001110001111010111000,
    22'b0001110100110011001101,
    22'b0001110100101000111101,
    22'b0001110110000101001000,
    22'b0001111000110011001101,
    22'b0001111001110000101001,
    22'b0001111000010100011111,
    22'b0001110110011001100110,
    22'b0001110100000000000000,
    22'b0001110011000010100100,
    22'b0001110010111000010100,
    22'b0001110010100011110110,
    22'b0001110010000101001000,
    22'b0001110001110000101001,
    22'b0001110001100110011010,
    22'b0001110001011100001010,
    22'b0001110000110011001101,
    22'b0001110000001010001111,
    22'b0001101111010111000011,
    22'b0001101111100001010010,
    22'b0001110000010100011111,
    22'b0001110000111101011100,
    22'b0001110000110011001101,
    22'b0001110000011110101110,
    22'b0001101111110101110001,
    22'b0001101101010001111011,
    22'b0001101010000101001000,
    22'b0001100110111000010100,
    22'b0001100100000000000000,
    22'b0001100001010001111011,
    22'b0001011101100110011010,
    22'b0001011001110000101001,
    22'b0001010111100001010010,
    22'b0001010101011100001010,
    22'b0001010011010111000011,
    22'b0001010001111010111000,
    22'b0001010001011100001010,
    22'b0001010001100110011010,
    22'b0001010001100110011010,
    22'b0001010010000101001000,
    22'b0001010100000000000000,
    22'b0001010110000101001000,
    22'b0001011000011110101110,
    22'b0001011011001100110011,
    22'b0001011111101011100001,
    22'b0001100010011001100110,
    22'b0001100100110011001101,
    22'b0001100110111000010100,
    22'b0001101000110011001101,
    22'b0001101001100110011010,
    22'b0001101001111010111000,
    22'b0001101001111010111000,
    22'b0001101001000111101100,
    22'b0001100101010001111011,
    22'b0001011110111000010100,
    22'b0001011011110101110001,
    22'b0001011011001100110011,
    22'b0001011011110101110001,
    22'b0001011011110101110001,
    22'b0001011000010100011111,
    22'b0001010100111101011100,
    22'b0001010010101110000101,
    22'b0001010000110011001101,
    22'b0001001101100110011010,
    22'b0001001011100001010010,
    22'b0001001000110011001101,
    22'b0001000110000101001000,
    22'b0000110011010111000011,
    22'b0000001011000010100100,
    22'b0000000010000101001000,
    22'b0000000000001010001111,
    22'b0000000000110011001101,
    22'b0000000011001100110011,
    22'b0000000110000101001000,
    22'b0000001010111000010100,
    22'b0000001011001100110011,
    22'b0000000111100001010010,
    22'b0000000011101011100001,
    22'b1111111100110011001101,
    22'b1111111001100110011010,
    22'b1111110110111000010100,
    22'b1111110010100011110110,
    22'b1111110001000111101100,
    22'b1111110001011100001010,
    22'b1111110010000101001000,
    22'b1111110011001100110011,
    22'b1111110101011100001010,
    22'b1111110101110000101001,
    22'b1111110101010001111011,
    22'b1111110100011110101110,
    22'b1111110100000000000000,
    22'b1111110010101110000101,
    22'b1111110010000101001000,
    22'b1111110010011001100110,
    22'b1111110100001010001111,
    22'b1111111000111101011100,
    22'b1111111101000111101100,
    22'b0000000001010001111011,
    22'b0000000101010001111011,
    22'b0000001000110011001101,
    22'b0000001100010100011111,
    22'b0000001110001111010111,
    22'b0000001111101011100001,
    22'b0000010001100110011010,
    22'b0000010101010001111011,
    22'b0000011111000010100100,
    22'b0000100101100110011010,
    22'b0000101011100001010010,
    22'b0000101111100001010010,
    22'b0000110000110011001101,
    22'b0000101111001100110011,
    22'b0000101101011100001010,
    22'b0000101010011001100110,
    22'b0000100111100001010010,
    22'b0000100100110011001101,
    22'b0000100010011001100110,
    22'b0000100001010001111011,
    22'b0000100000000000000000,
    22'b0000011110101110000101,
    22'b0000011101011100001010,
    22'b0000011100010100011111,
    22'b0000011011110101110001,
    22'b0000011100000000000000,
    22'b0000011100011110101110,
    22'b0000011101011100001010,
    22'b0000011110011001100110,
    22'b0000011110011001100110,
    22'b0000011101110000101001,
    22'b0000011100101000111101,
    22'b0000011011000010100100,
    22'b0000011001011100001010,
    22'b0000011000001010001111,
    22'b0000010111101011100001,
    22'b0000010111010111000011,
    22'b0000011000000000000000,
    22'b0000011001100110011010,
    22'b0000011011110101110001,
    22'b0000011110011001100110,
    22'b0000100000111101011100,
    22'b0000100011010111000011,
    22'b0000100110100011110110,
    22'b0000101001010001111011,
    22'b0000101100011110101110,
    22'b0000101111010111000011,
    22'b0000110010001111010111,
    22'b0000110111000010100100,
    22'b0000111001111010111000,
    22'b0000111011000010100100,
    22'b0000111011110101110001,
    22'b0000111100010100011111,
    22'b0000111100011110101110,
    22'b0000111010000101001000,
    22'b0000111000001010001111,
    22'b0000110110101110000101,
    22'b0000110101011100001010,
    22'b0000110010101110000101,
    22'b0000110001110000101001,
    22'b0000110000101000111101,
    22'b0000101111001100110011,
    22'b0000101100000000000000,
    22'b0000101001111010111000,
    22'b0000100110011001100110,
    22'b0000100100001010001111,
    22'b0000100001100110011010,
    22'b0000100100011110101110,
    22'b0000100111110101110001,
    22'b0000101100111101011100,
    22'b0000110000111101011100,
    22'b0000110101010001111011,
    22'b0000111110011001100110,
    22'b0001000110001111010111,
    22'b0001001101011100001010,
    22'b0001001101111010111000,
    22'b0001001000101000111101,
    22'b0001000000010100011111,
    22'b0000111011000010100100,
    22'b0000110110001111010111,
    22'b0000110010001111010111,
    22'b0000101111010111000011,
    22'b0000101111100001010010,
    22'b0000110000101000111101,
    22'b0000110010001111010111,
    22'b0000110011101011100001,
    22'b0000110100111101011100,
    22'b0000110100110011001101,
    22'b0000110011100001010010,
    22'b0000110001110000101001,
    22'b0000101111010111000011,
    22'b0000101101110000101001,
    22'b0000101100010100011111,
    22'b0000101010111000010100,
    22'b0000101001011100001010,
    22'b0000100111010111000011,
    22'b0000100100111101011100,
    22'b0000100011001100110011,
    22'b0000100000010100011111,
    22'b0000011110011001100110,
    22'b0000011110011001100110,
    22'b0000011101111010111000,
    22'b0000011110001111010111,
    22'b0000011110001111010111,
    22'b0000011111110101110001,
    22'b0000100000001010001111,
    22'b0000100001110000101001,
    22'b0000100100000000000000,
    22'b0000100110011001100110,
    22'b0000101010000101001000,
    22'b0000101100010100011111,
    22'b0000101101011100001010,
    22'b0000101111001100110011,
    22'b0000101111001100110011,
    22'b0000101101100110011010,
    22'b0000101100011110101110,
    22'b0000101011000010100100,
    22'b0000101001111010111000,
    22'b0000101000001010001111,
    22'b0000100100111101011100,
    22'b0000100010000101001000,
    22'b0000011110100011110110,
    22'b0000011001100110011010,
    22'b0000010101010001111011,
    22'b0000010000110011001101,
    22'b0000001100110011001101,
    22'b0000001010001111010111,
    22'b0000001000101000111101,
    22'b0000001000110011001101,
    22'b0000001010000101001000,
    22'b0000001011000010100100,
    22'b0000001100010100011111,
    22'b0000001110101110000101,
    22'b0000010010011001100110,
    22'b0000010101010001111011,
    22'b0000010111001100110011,
    22'b0000010100010100011111,
    22'b0000010110000101001000,
    22'b0000011100101000111101,
    22'b0000100011110101110001,
    22'b0000101001100110011010,
    22'b0000101101010001111011,
    22'b0000101011100001010010,
    22'b0000101101000111101100,
    22'b0000110001010001111011,
    22'b0000110101010001111011,
    22'b0000111001000111101100,
    22'b0000111100011110101110,
    22'b0000111011101011100001,
    22'b0000111001100110011010,
    22'b0000110111110101110001,
    22'b0000110011010111000011,
    22'b0000101100000000000000,
    22'b0000100101011100001010,
    22'b0000100001000111101100,
    22'b0000011111100001010010,
    22'b0000100000110011001101,
    22'b0000100100001010001111,
    22'b0000100111001100110011,
    22'b0000101000110011001101,
    22'b0000101010001111010111,
    22'b0000101111000010100100,
    22'b0000101101011100001010,
    22'b0000101001110000101001,
    22'b0000100100111101011100,
    22'b0000011100000000000000,
    22'b0000010110001111010111,
    22'b0000010000101000111101,
    22'b0000001011100001010010,
    22'b0000000101111010111000,
    22'b1111111101011100001010,
    22'b1111110111101011100001,
    22'b1111110011100001010010,
    22'b1111110000011110101110,
    22'b1111101101111010111000,
    22'b1111101101000111101100,
    22'b1111101100110011001101,
    22'b1111101100110011001101,
    22'b1111101101000111101100,
    22'b1111101101011100001010,
    22'b1111101110000101001000,
    22'b1111101111001100110011,
    22'b1111110000101000111101,
    22'b1111110011001100110011,
    22'b1111110101011100001010,
    22'b1111110111101011100001,
    22'b1111111001111010111000,
    22'b1111111100011110101110,
    22'b1111111110011001100110,
    22'b1111111111110101110001,
    22'b0000000001010001111011,
    22'b0000000010101110000101,
    22'b0000000100001010001111,
    22'b0000000101010001111011,
    22'b0000000100010100011111,
    22'b0000000111100001010010,
    22'b0000001010001111010111,
    22'b0000001011100001010010,
    22'b0000001101000111101100,
    22'b0000001110100011110110,
    22'b0000010000010100011111,
    22'b0000010100010100011111,
    22'b0000010110001111010111,
    22'b0000010111101011100001,
    22'b0000011001011100001010,
    22'b0000011000011110101110,
    22'b0000011001010001111011,
    22'b0000010011000010100100,
    22'b0000001000001010001111,
    22'b1111111011101011100001,
    22'b1111100111001100110011,
    22'b1111011101011100001010,
    22'b1111100100011110101110,
    22'b1111110111110101110001,
    22'b1111111101111010111000,
    22'b1111111101010001111011,
    22'b0000001010000101001000,
    22'b0000011111010111000011,
    22'b0000100100101000111101,
    22'b0000100011010111000011,
    22'b0000100000000000000000,
    22'b0000011110100011110110,
    22'b0000010110001111010111,
    22'b0000001111110101110001,
    22'b0000001100110011001101,
    22'b0000001101010001111011,
    22'b0000001111000010100100,
    22'b0000010001111010111000,
    22'b0000010100010100011111,
    22'b0000010110101110000101,
    22'b0000011001010001111011,
    22'b0000011101110000101001,
    22'b0000100001011100001010,
    22'b0000100100110011001101,
    22'b0000100111101011100001,
    22'b0000101001110000101001,
    22'b0000101011001100110011,
    22'b0000101010101110000101,
    22'b0000101000110011001101,
    22'b0000100101110000101001,
    22'b0000100001100110011010,
    22'b0000011110000101001000,
    22'b0000011001111010111000,
    22'b0000010101000111101100,
    22'b0000001101110000101001,
    22'b0000001001010001111011,
    22'b0000000101010001111011,
    22'b0000000001000111101100,
    22'b1111111100111101011100,
    22'b1111111011000010100100,
    22'b1111111001100110011010,
    22'b1111110111010111000011,
    22'b1111110100111101011100,
    22'b1111110011101011100001,
    22'b1111110010101110000101,
    22'b1111110000110011001101,
    22'b1111101111110101110001,
    22'b1111110000001010001111,
    22'b1111110000110011001101,
    22'b1111110001011100001010,
    22'b1111110001111010111000,
    22'b1111110001010001111011,
    22'b1111110001111010111000,
    22'b1111110010100011110110,
    22'b1111110011000010100100,
    22'b1111110011100001010010,
    22'b1111110011110101110001,
    22'b1111110100010100011111,
    22'b1111110100111101011100,
    22'b1111110101100110011010,
    22'b1111110110101110000101,
    22'b1111110111100001010010,
    22'b1111111000011110101110,
    22'b1111111001010001111011,
    22'b1111111010100011110110,
    22'b1111111011010111000011,
    22'b1111111100000000000000,
    22'b1111111100110011001101,
    22'b1111111101110000101001,
    22'b1111111110100011110110,
    22'b1111111111010111000011,
    22'b0000000000001010001111,
    22'b0000000001000111101100,
    22'b0000000010100011110110,
    22'b0000000011101011100001,
    22'b0000000101000111101100,
    22'b0000000110100011110110,
    22'b0000000111101011100001,
    22'b0000001001010001111011,
    22'b0000001010001111010111,
    22'b0000001011000010100100,
    22'b0000001011010111000011,
    22'b0000001011101011100001,
    22'b0000001011101011100001,
    22'b0000001011001100110011,
    22'b0000001010100011110110,
    22'b0000001010000101001000,
    22'b0000001001100110011010,
    22'b0000001000110011001101,
    22'b0000000111110101110001,
    22'b0000000110111000010100,
    22'b0000000101110000101001,
    22'b0000000100110011001101,
    22'b0000000011110101110001,
    22'b0000000011010111000011,
    22'b0000000010101110000101,
    22'b0000000010001111010111,
    22'b0000000001100110011010,
    22'b0000000000111101011100,
    22'b0000000000010100011111,
    22'b0000000000010100011111,
    22'b0000000000000000000000,
    22'b1111111111101011100001,
    22'b1111111110011001100110,
    22'b1111111110001111010111,
    22'b1111111101110000101001,
    22'b1111111101010001111011,
    22'b1111111100001010001111,
    22'b1111110101010001111011,
    22'b1111110011101011100001,
    22'b1111110101000111101100,
    22'b1111110110111000010100,
    22'b1111110101100110011010,
    22'b1111110101000111101100,
    22'b1111110101010001111011,
    22'b1111110110001111010111,
    22'b1111111000000000000000,
    22'b1111111000111101011100,
    22'b1111111001100110011010,
    22'b1111111010001111010111,
    22'b1111111010100011110110,
    22'b1111111010100011110110,
    22'b1111111010011001100110,
    22'b1111111010001111010111,
    22'b1111111001111010111000,
    22'b1111111001011100001010,
    22'b1111111001000111101100,
    22'b1111111000110011001101,
    22'b1111111000101000111101,
    22'b1111111000011110101110,
    22'b1111111000011110101110,
    22'b1111111000101000111101,
    22'b1111111000101000111101,
    22'b1111111000110011001101,
    22'b1111111000110011001101,
    22'b1111111000110011001101,
    22'b1111111000101000111101,
    22'b1111111000010100011111,
    22'b1111111000000000000000,
    22'b1111110111100001010010,
    22'b1111110111001100110011,
    22'b1111110110101110000101,
    22'b1111110110011001100110,
    22'b1111110110000101001000,
    22'b1111110101111010111000,
    22'b1111110101110000101001,
    22'b1111110101011100001010,
    22'b1111110101010001111011,
    22'b1111110101000111101100,
    22'b1111110100111101011100,
    22'b1111110100110011001101,
    22'b1111110100101000111101,
    22'b1111110100011110101110,
    22'b1111110100001010001111,
    22'b1111110011101011100001,
    22'b1111110011000010100100,
    22'b1111110010011001100110,
    22'b1111110001100110011010,
    22'b1111110001000111101100,
    22'b1111110000111101011100,
    22'b1111110000101000111101,
    22'b1111101111110101110001,
    22'b1111101111000010100100,
    22'b1111101011100001010010,
    22'b1111100110101110000101,
    22'b1111100110011001100110,
    22'b1111100111110101110001,
    22'b1111101001100110011010,
    22'b1111101011100001010010,
    22'b1111101101110000101001,
    22'b1111101111010111000011,
    22'b1111110001000111101100,
    22'b1111110011010111000011,
    22'b1111110110101110000101,
    22'b1111111001011100001010,
    22'b1111111100011110101110,
    22'b0000000000011110101110,
    22'b0000000011100001010010,
    22'b0000000110100011110110,
    22'b0000001001110000101001,
    22'b0000001100110011001101,
    22'b0000010000010100011111,
    22'b0000010010100011110110,
    22'b0000010100101000111101,
    22'b0000010110011001100110,
    22'b0000011000011110101110,
    22'b0000011001100110011010,
    22'b0000011001111010111000,
    22'b0000011001100110011010,
    22'b0000011000110011001101,
    22'b0000010111110101110001,
    22'b0000010110011001100110,
    22'b0000010100001010001111,
    22'b0000001110101110000101,
    22'b0000001011100001010010,
    22'b0000000110100011110110,
    22'b0000000100111101011100,
    22'b0000000011110101110001,
    22'b0000000010000101001000,
    22'b0000000000110011001101,
    22'b0000000000001010001111,
    22'b1111111111000010100100,
    22'b1111111110000101001000,
    22'b1111111110000101001000,
    22'b1111111110100011110110,
    22'b0000001011000010100100,
    22'b0000001101000111101100,
    22'b0000001110100011110110,
    22'b0000001110111000010100,
    22'b0000001110111000010100,
    22'b0000001110001111010111,
    22'b0000001100101000111101,
    22'b0000001011101011100001,
    22'b0000001010001111010111,
    22'b0000001000110011001101,
    22'b0000000111000010100100,
    22'b0000000110100011110110,
    22'b0000000101111010111000,
    22'b0000000101110000101001,
    22'b0000000101100110011010,
    22'b0000000101010001111011,
    22'b0000000100110011001101,
    22'b0000000100011110101110,
    22'b0000000100001010001111,
    22'b0000000100001010001111,
    22'b0000000100101000111101,
    22'b0000000101100110011010,
    22'b0000000111110101110001,
    22'b0000001001100110011010,
    22'b0000001011101011100001,
    22'b0000001110000101001000,
    22'b0000001111110101110001,
    22'b0000010001010001111011,
    22'b0000010010100011110110,
    22'b0000010100000000000000,
    22'b0000010100111101011100,
    22'b0000010101111010111000,
    22'b0000010110111000010100,
    22'b0000010111110101110001,
    22'b0000010110001111010111,
    22'b0000010110100011110110,
    22'b0000010111001100110011,
    22'b0000010110111000010100,
    22'b0000010110101110000101,
    22'b0000010110100011110110,
    22'b0000010111101011100001,
    22'b0000011000000000000000,
    22'b0000011000110011001101,
    22'b0000011100000000000000,
    22'b0000100000010100011111,
    22'b0000100100011110101110,
    22'b0000100111110101110001,
    22'b0000101010011001100110,
    22'b0000101100000000000000,
    22'b0000101010011001100110,
    22'b0000101000110011001101,
    22'b0000100110011001100110,
    22'b0000100010000101001000,
    22'b0000011101111010111000,
    22'b0000011000111101011100,
    22'b0000010101100110011010,
    22'b0000010000110011001101,
    22'b0000000101011100001010,
    22'b0000000011001100110011,
    22'b1111111111101011100001,
    22'b1111111100111101011100,
    22'b1111111010011001100110,
    22'b1111111000001010001111,
    22'b1111110110001111010111,
    22'b1111110101011100001010,
    22'b1111110100111101011100,
    22'b1111110100010100011111,
    22'b1111110100000000000000,
    22'b1111110011101011100001,
    22'b1111110011100001010010,
    22'b1111110011100001010010,
    22'b1111110011100001010010,
    22'b1111110011101011100001,
    22'b1111110011110101110001,
    22'b1111110011110101110001,
    22'b1111110011010111000011,
    22'b1111110010001111010111,
    22'b1111101111110101110001,
    22'b1111101101011100001010,
    22'b1111101011000010100100,
    22'b1111101000101000111101,
    22'b1111100110011001100110,
    22'b1111100110000101001000,
    22'b1111100111001100110011,
    22'b1111101001110000101001,
    22'b1111101101000111101100,
    22'b1111101111010111000011,
    22'b1111110001000111101100,
    22'b1111110011001100110011,
    22'b1111110100111101011100,
    22'b1111110110101110000101,
    22'b1111111000011110101110,
    22'b1111111010011001100110,
    22'b1111111011001100110011,
    22'b1111111011010111000011,
    22'b1111111010011001100110,
    22'b1111111000110011001101,
    22'b1111110010111000010100,
    22'b1111110010100011110110,
    22'b1111110010011001100110,
    22'b1111110010001111010111,
    22'b1111110010001111010111,
    22'b1111110001111010111000,
    22'b1111110001100110011010,
    22'b1111110000111101011100,
    22'b1111110000010100011111,
    22'b1111101111010111000011,
    22'b1111101110111000010100,
    22'b1111101111000010100100,
    22'b1111101110101110000101,
    22'b1111101110000101001000,
    22'b1111101101100110011010,
    22'b1111101101000111101100,
    22'b1111101100101000111101,
    22'b1111101100011110101110,
    22'b1111101100011110101110,
    22'b1111101100101000111101,
    22'b1111101100010100011111,
    22'b1111101011110101110001,
    22'b1111101011001100110011,
    22'b1111101010001111010111,
    22'b1111101001010001111011,
    22'b1111101000011110101110,
    22'b1111100111010111000011,
    22'b1111100101110000101001,
    22'b1111100100011110101110,
    22'b1111100011000010100100,
    22'b1111100001100110011010,
    22'b1111100000000000000000,
    22'b1111010110000101001000,
    22'b1111010100010100011111,
    22'b1111010010101110000101,
    22'b1111010001011100001010,
    22'b1111001111110101110001,
    22'b1111001101111010111000,
    22'b1111001011110101110001,
    22'b1111001001111010111000,
    22'b1111001000111101011100,
    22'b1111001011100001010010,
    22'b1111001101110000101001,
    22'b1111010001111010111000,
    22'b1111010100111101011100,
    22'b1111010101110000101001,
    22'b1111010101111010111000,
    22'b1111010111100001010010,
    22'b1111011011101011100001,
    22'b1111011111010111000011,
    22'b1111100000101000111101,
    22'b1111011110111000010100,
    22'b1111011000011110101110,
    22'b1111010101000111101100,
    22'b1111010001000111101100,
    22'b1111001110111000010100,
    22'b1111001110001111010111,
    22'b1111001101100110011010,
    22'b1111001101110000101001,
    22'b1111001110101110000101,
    22'b1111001111000010100100,
    22'b1111001111100001010010,
    22'b1111010000110011001101,
    22'b1111010101010001111011,
    22'b1111011001111010111000,
    22'b1111011101111010111000,
    22'b1111101000110011001101,
    22'b1111101010100011110110,
    22'b1111101100001010001111,
    22'b1111101101111010111000,
    22'b1111101111100001010010,
    22'b1111101111110101110001,
    22'b1111101111100001010010,
    22'b1111101111000010100100,
    22'b1111101101111010111000,
    22'b1111101101010001111011,
    22'b1111101100110011001101,
    22'b1111101100101000111101,
    22'b1111101100011110101110,
    22'b1111101100010100011111,
    22'b1111101100011110101110,
    22'b1111101100101000111101,
    22'b1111101100010100011111,
    22'b1111101100001010001111,
    22'b1111101100010100011111,
    22'b1111101100101000111101,
    22'b1111101100110011001101,
    22'b1111101101000111101100,
    22'b1111101101000111101100,
    22'b1111101100110011001101,
    22'b1111101100010100011111,
    22'b1111101011110101110001,
    22'b1111101011010111000011,
    22'b1111101010101110000101,
    22'b1111101010100011110110,
    22'b1111101010111000010100,
    22'b1111101011000010100100,
    22'b1111101011110101110001,
    22'b1111101100000000000000,
    22'b1111101011110101110001,
    22'b1111101011110101110001,
    22'b1111101100000000000000,
    22'b1111101011110101110001,
    22'b1111101100010100011111,
    22'b1111101101110000101001,
    22'b1111101111010111000011,
    22'b1111110000010100011111,
    22'b1111110001000111101100,
    22'b1111110001110000101001,
    22'b1111110001110000101001,
    22'b1111110001100110011010,
    22'b1111110010011001100110,
    22'b1111110011001100110011,
    22'b1111110011110101110001,
    22'b1111110101100110011010,
    22'b1111111000011110101110,
    22'b1111111011100001010010,
    22'b1111111110101110000101,
    22'b0000000001011100001010,
    22'b0000000100011110101110,
    22'b0000000110011001100110,
    22'b0000000111010111000011,
    22'b0000001011001100110011,
    22'b0000001100101000111101,
    22'b0000001101100110011010,
    22'b0000001110101110000101,
    22'b0000001101110000101001,
    22'b0000001001111010111000,
    22'b0000000110100011110110,
    22'b0000000011000010100100,
    22'b1111111110111000010100,
    22'b1111111101010001111011,
    22'b1111111100001010001111,
    22'b1111111011100001010010,
    22'b1111111011010111000011,
    22'b1111111011010111000011,
    22'b1111111011110101110001,
    22'b1111111100010100011111,
    22'b1111111100101000111101,
    22'b1111111110000101001000,
    22'b0000000000000000000000,
    22'b0000000001100110011010,
    22'b0000000011000010100100,
    22'b0000000100111101011100,
    22'b0000000111101011100001,
    22'b0000001001000111101100,
    22'b0000001001110000101001,
    22'b0000001010111000010100,
    22'b0000001100010100011111,
    22'b0000001101100110011010,
    22'b0000001110101110000101,
    22'b0000010000001010001111,
    22'b0000001111000010100100,
    22'b0000001011010111000011,
    22'b0000000111110101110001,
    22'b0000000101111010111000,
    22'b0000000100101000111101,
    22'b0000000011010111000011,
    22'b0000000001110000101001,
    22'b0000000000101000111101,
    22'b1111111111001100110011,
    22'b1111111101111010111000,
    22'b1111111100010100011111,
    22'b1111111011000010100100,
    22'b1111111001111010111000,
    22'b1111111000111101011100,
    22'b1111111000010100011111,
    22'b1111111000110011001101,
    22'b1111111001010001111011,
    22'b1111111001110000101001,
    22'b1111111010001111010111,
    22'b1111111010111000010100,
    22'b1111111011101011100001,
    22'b1111111100010100011111,
    22'b1111111101110000101001,
    22'b1111111111101011100001,
    22'b0000000001000111101100,
    22'b0000000011100001010010,
    22'b0000000110000101001000,
    22'b0000000111101011100001,
    22'b0000000111000010100100,
    22'b0000001001111010111000,
    22'b0000010001000111101100,
    22'b0000011000011110101110,
    22'b0000100001010001111011,
    22'b0000100100101000111101,
    22'b0000100100000000000000,
    22'b0000100001011100001010,
    22'b0000011110101110000101,
    22'b0000011011101011100001,
    22'b0000011000000000000000,
    22'b0000010101110000101001,
    22'b0000010100011110101110,
    22'b0000010011100001010010,
    22'b0000010010001111010111,
    22'b0000010001100110011010,
    22'b0000010001011100001010,
    22'b0000010001100110011010,
    22'b0000010001100110011010,
    22'b0000010001010001111011,
    22'b0000010000110011001101,
    22'b0000010000001010001111,
    22'b0000001111100001010010,
    22'b0000001110001111010111,
    22'b0000001101010001111011,
    22'b0000001011110101110001,
    22'b0000001010100011110110,
    22'b0000001001000111101100,
    22'b0000001000111101011100,
    22'b0000001001010001111011,
    22'b0000001001110000101001,
    22'b0000001010001111010111,
    22'b0000001010101110000101,
    22'b0000001011001100110011,
    22'b0000001011110101110001,
    22'b0000001101011100001010,
    22'b0000001111100001010010,
    22'b0000010001000111101100,
    22'b0000010001111010111000,
    22'b0000010010000101001000,
    22'b0000010000110011001101,
    22'b0000001110011001100110,
    22'b0000001011000010100100,
    22'b0000001000110011001101,
    22'b0000000110100011110110,
    22'b0000000100011110101110,
    22'b0000000010101110000101,
    22'b0000000001110000101001,
    22'b0000000001000111101100,
    22'b0000000000011110101110,
    22'b0000000000000000000000,
    22'b1111111111110101110001,
    22'b1111111111000010100100,
    22'b1111111111000010100100,
    22'b1111111110001111010111,
    22'b1111111100101000111101,
    22'b1111111010111000010100,
    22'b1111111000111101011100,
    22'b1111110110011001100110,
    22'b1111110100110011001101,
    22'b1111110011001100110011,
    22'b1111110010000101001000,
    22'b1111110001000111101100,
    22'b1111110000110011001101,
    22'b1111110000110011001101,
    22'b1111110001000111101100,
    22'b1111110001110000101001,
    22'b1111110010000101001000,
    22'b1111110001000111101100,
    22'b1111101111010111000011,
    22'b1111101110011001100110,
    22'b1111101101100110011010,
    22'b1111101011000010100100,
    22'b1111101000000000000000,
    22'b1111100111010111000011,
    22'b1111101001111010111000,
    22'b1111100100110011001101,
    22'b1111100111000010100100,
    22'b1111100111101011100001,
    22'b1111100111110101110001,
    22'b1111100111110101110001,
    22'b1111101000111101011100,
    22'b1111101001010001111011,
    22'b1111100111010111000011,
    22'b1111101000110011001101,
    22'b1111101011010111000011,
    22'b1111101100101000111101,
    22'b1111101011001100110011,
    22'b1111101000000000000000,
    22'b1111100111110101110001,
    22'b1111100111101011100001,
    22'b1111100111001100110011,
    22'b1111100111100001010010,
    22'b1111101000111101011100,
    22'b1111101001010001111011,
    22'b1111101001110000101001,
    22'b1111101011001100110011,
    22'b1111101100110011001101,
    22'b1111101110011001100110,
    22'b1111110000001010001111,
    22'b1111110001011100001010,
    22'b1111110010011001100110,
    22'b1111110101000111101100,
    22'b1111110100010100011111,
    22'b1111110010101110000101,
    22'b1111110000110011001101,
    22'b1111101110000101001000,
    22'b1111101100001010001111,
    22'b1111101010001111010111,
    22'b1111101000111101011100,
    22'b1111101000011110101110,
    22'b1111101000001010001111,
    22'b1111101000000000000000,
    22'b1111101010000101001000,
    22'b1111101011101011100001,
    22'b1111101101000111101100,
    22'b1111101110101110000101,
    22'b1111110000000000000000,
    22'b1111110000101000111101,
    22'b1111110001010001111011,
    22'b1111110001110000101001,
    22'b1111110001111010111000,
    22'b1111110001100110011010,
    22'b1111110001010001111011,
    22'b1111110001010001111011,
    22'b1111110001011100001010,
    22'b1111110001010001111011,
    22'b1111110000111101011100,
    22'b1111101111110101110001,
    22'b1111101110101110000101,
    22'b1111101110011001100110,
    22'b1111101110011001100110,
    22'b1111101110100011110110,
    22'b1111101110100011110110,
    22'b1111101101111010111000,
    22'b1111101101010001111011,
    22'b1111101101011100001010,
    22'b1111101101111010111000,
    22'b1111101110100011110110,
    22'b1111101111100001010010,
    22'b1111110001010001111011,
    22'b1111110010100011110110,
    22'b1111110011101011100001,
    22'b1111110100011110101110,
    22'b1111110100011110101110,
    22'b1111110100011110101110,
    22'b1111110100101000111101,
    22'b1111110101000111101100,
    22'b1111110101110000101001,
    22'b1111110110011001100110,
    22'b1111110111000010100100,
    22'b1111110111110101110001,
    22'b1111111001010001111011,
    22'b1111111010011001100110,
    22'b1111111011000010100100,
    22'b1111111011110101110001,
    22'b1111111100110011001101,
    22'b1111111101100110011010,
    22'b1111111101100110011010,
    22'b1111111101100110011010,
    22'b1111111101011100001010,
    22'b1111111101000111101100,
    22'b1111111101000111101100,
    22'b1111111101000111101100,
    22'b1111111100111101011100,
    22'b1111111100011110101110,
    22'b1111111011110101110001,
    22'b1111111011010111000011,
    22'b1111111010101110000101,
    22'b1111111010001111010111,
    22'b1111111010000101001000,
    22'b1111111010001111010111,
    22'b1111111010101110000101,
    22'b1111111011010111000011,
    22'b1111111100000000000000,
    22'b1111101111100001010010,
    22'b1111101011100001010010,
    22'b1111101000001010001111,
    22'b1111100011100001010010,
    22'b1111100001111010111000,
    22'b1111100010011001100110,
    22'b1111100001000111101100,
    22'b1111011111000010100100,
    22'b1111011111101011100001,
    22'b1111011111101011100001,
    22'b1111100000010100011111,
    22'b1111100010101110000101,
    22'b1111100100111101011100,
    22'b1111100111010111000011,
    22'b1111101010111000010100,
    22'b1111101110001111010111,
    22'b1111110010000101001000,
    22'b1111110100010100011111,
    22'b1111110110000101001000,
    22'b1111110111000010100100,
    22'b1111110111101011100001,
    22'b1111110111101011100001,
    22'b1111110111001100110011,
    22'b1111110110111000010100,
    22'b1111110110101110000101,
    22'b1111110110011001100110,
    22'b1111110110011001100110,
    22'b1111110110101110000101,
    22'b1111110111000010100100,
    22'b1111110110111000010100,
    22'b1111110111000010100100,
    22'b1111110111001100110011,
    22'b1111110110101110000101,
    22'b1111110110011001100110,
    22'b1111110111000010100100,
    22'b1111110111110101110001,
    22'b1111111000110011001101,
    22'b1111111001110000101001,
    22'b1111111011001100110011,
    22'b1111111100110011001101,
    22'b1111111110101110000101,
    22'b0000000000001010001111,
    22'b0000000001011100001010,
    22'b0000000010011001100110,
    22'b0000000011000010100100,
    22'b0000000011001100110011,
    22'b0000000011001100110011,
    22'b0000000011010111000011,
    22'b0000000011100001010010,
    22'b0000000011001100110011,
    22'b0000000011000010100100,
    22'b0000000010101110000101,
    22'b0000000010101110000101,
    22'b0000000011000010100100,
    22'b0000000011001100110011,
    22'b0000000010111000010100,
    22'b0000000001111010111000,
    22'b0000000010001111010111,
    22'b0000000010000101001000,
    22'b0000001010000101001000,
    22'b0000001011000010100100,
    22'b0000001100011110101110,
    22'b0000001110000101001000,
    22'b0000010000000000000000,
    22'b0000010001000111101100,
    22'b0000010010000101001000,
    22'b0000010010100011110110,
    22'b0000010011000010100100,
    22'b0000010011001100110011,
    22'b0000010011010111000011,
    22'b0000010011100001010010,
    22'b0000010011101011100001,
    22'b0000010100010100011111,
    22'b0000010100011110101110,
    22'b0000010100111101011100,
    22'b0000010101110000101001,
    22'b0000010111001100110011,
    22'b0000011000010100011111,
    22'b0000011001100110011010,
    22'b0000011010101110000101,
    22'b0000011100001010001111,
    22'b0000011101000111101100,
    22'b0000011101110000101001,
    22'b0000011110100011110110,
    22'b0000011110111000010100,
    22'b0000011111000010100100,
    22'b0000011111001100110011,
    22'b0000011111000010100100,
    22'b0000011110111000010100,
    22'b0000011110011001100110,
    22'b0000011101110000101001,
    22'b0000011100011110101110,
    22'b0000011011001100110011,
    22'b0000011001110000101001,
    22'b0000011000001010001111,
    22'b0000010110001111010111,
    22'b0000010100110011001101,
    22'b0000010011100001010010,
    22'b0000010010000101001000,
    22'b0000010000011110101110,
    22'b0000001111001100110011,
    22'b0000001101111010111000,
    22'b0000001100101000111101,
    22'b0000001010111000010100,
    22'b0000001001100110011010,
    22'b0000001000011110101110,
    22'b0000000111100001010010,
    22'b0000000010001111010111,
    22'b0000000000110011001101,
    22'b1111111111100001010010,
    22'b1111111100111101011100,
    22'b1111111010001111010111,
    22'b1111110111101011100001,
    22'b1111110100011110101110,
    22'b1111101110100011110110,
    22'b1111101010001111010111,
    22'b1111100001111010111000,
    22'b1111011000011110101110,
    22'b1111101000001010001111,
    22'b1111110100110011001101,
    22'b1111110101011100001010,
    22'b0000000000110011001101,
    22'b0000000011100001010010,
    22'b1111111011010111000011,
    22'b1111110110011001100110,
    22'b1111110010011001100110,
    22'b1111101110001111010111,
    22'b1111101111110101110001,
    22'b1111110010101110000101,
    22'b1111110011010111000011,
    22'b1111110010000101001000,
    22'b1111101111100001010010,
    22'b1111101100000000000000,
    22'b1111100111100001010010,
    22'b1111100101011100001010,
    22'b1111100100001010001111,
    22'b1111100100000000000000,
    22'b1111100100101000111101,
    22'b1111100101011100001010,
    22'b1111100110000101001000,
    22'b1111100110100011110110,
    22'b1111100110001111010111,
    22'b1111100101011100001010,
    22'b1111100100011110101110,
    22'b1111100011110101110001,
    22'b1111100011110101110001,
    22'b1111100011010111000011,
    22'b1111100010101110000101,
    22'b1111100001100110011010,
    22'b1111100000110011001101,
    22'b1111100000010100011111,
    22'b1111100000010100011111,
    22'b1111100000000000000000,
    22'b1111011111110101110001,
    22'b1111100000000000000000,
    22'b1111011111110101110001,
    22'b1111011111110101110001,
    22'b1111100000000000000000,
    22'b1111100000001010001111,
    22'b1111100000101000111101,
    22'b1111100001010001111011,
    22'b1111100001110000101001,
    22'b1111100010001111010111,
    22'b1111100010111000010100,
    22'b1111100011000010100100,
    22'b1111100011010111000011,
    22'b1111100011100001010010,
    22'b1111100011101011100001,
    22'b1111100100001010001111,
    22'b1111100100001010001111,
    22'b1111100100000000000000,
    22'b1111100100001010001111,
    22'b1111100101010001111011,
    22'b1111100101111010111000,
    22'b1111100110111000010100,
    22'b1111101001000111101100,
    22'b1111101010011001100110,
    22'b1111101011010111000011,
    22'b1111101100010100011111,
    22'b1111101100111101011100,
    22'b1111101101100110011010,
    22'b1111101110011001100110,
    22'b1111101111001100110011,
    22'b1111110000011110101110,
    22'b1111110100001010001111,
    22'b1111110101000111101100,
    22'b1111110110000101001000,
    22'b1111110110100011110110,
    22'b1111110110101110000101,
    22'b1111110110000101001000,
    22'b1111110100111101011100,
    22'b1111110101111010111000,
    22'b1111110111001100110011,
    22'b1111111000111101011100,
    22'b1111111010000101001000,
    22'b1111111011000010100100,
    22'b1111111100000000000000,
    22'b1111111101000111101100,
    22'b1111111101111010111000,
    22'b1111111111000010100100,
    22'b0000000000000000000000,
    22'b0000000000101000111101,
    22'b0000000001010001111011,
    22'b0000000001111010111000,
    22'b0000000010100011110110,
    22'b0000000011000010100100,
    22'b0000000011100001010010,
    22'b0000000100010100011111,
    22'b0000000100110011001101,
    22'b0000000100111101011100,
    22'b0000000101000111101100,
    22'b0000000100111101011100,
    22'b0000000100000000000000,
    22'b0000000001100110011010,
    22'b1111111111101011100001,
    22'b1111111101011100001010,
    22'b1111111010100011110110,
    22'b1111111001010001111011,
    22'b1111111001100110011010,
    22'b1111111010001111010111,
    22'b1111111010000101001000,
    22'b1111111001110000101001,
    22'b1111111001100110011010,
    22'b1111111001000111101100,
    22'b1111111001010001111011,
    22'b1111111010001111010111,
    22'b1111111011000010100100,
    22'b1111111011100001010010,
    22'b1111111100000000000000,
    22'b1111111100111101011100,
    22'b1111111100111101011100,
    22'b1111111100110011001101,
    22'b1111111101010001111011,
    22'b1111111101111010111000,
    22'b0000000000010100011111,
    22'b0000000010000101001000,
    22'b0000000011100001010010,
    22'b0000000101000111101100,
    22'b0000000110011001100110,
    22'b0000000101110000101001,
    22'b0000000101110000101001,
    22'b0000000101010001111011,
    22'b0000000100101000111101,
    22'b0000000011000010100100,
    22'b0000000010000101001000,
    22'b0000000000111101011100,
    22'b1111111111110101110001,
    22'b1111111110100011110110,
    22'b1111111110000101001000,
    22'b1111111110000101001000,
    22'b1111111101111010111000,
    22'b1111111110100011110110,
    22'b0000000000110011001101,
    22'b0000000011000010100100,
    22'b0000000101011100001010,
    22'b0000001000101000111101,
    22'b0000001011101011100001,
    22'b0000001110111000010100,
    22'b0000010001011100001010,
    22'b0000010100101000111101,
    22'b0000010111100001010010,
    22'b0000010111100001010010,
    22'b0000010101000111101100,
    22'b0000010010111000010100,
    22'b0000010000111101011100,
    22'b0000001111001100110011,
    22'b0000001100110011001101,
    22'b0000001010001111010111,
    22'b0000000111100001010010,
    22'b0000000100101000111101,
    22'b0000000010001111010111,
    22'b1111111111110101110001,
    22'b1111111110100011110110,
    22'b1111111101100110011010,
    22'b1111111100101000111101,
    22'b1111111100010100011111,
    22'b1111111100111101011100,
    22'b1111111110111000010100,
    22'b0000000101110000101001,
    22'b0000010101110000101001,
    22'b0000011100110011001101,
    22'b0000100010011001100110,
    22'b0000101101010001111011,
    22'b0000110101111010111000,
    22'b0000111011010111000011,
    22'b0000111100001010001111,
    22'b0000111000011110101110,
    22'b0000110011101011100001,
    22'b0000101101110000101001,
    22'b0000100111110101110001,
    22'b0000100001100110011010,
    22'b0000011011110101110001,
    22'b0000010101111010111000,
    22'b0000001110100011110110,
    22'b0000001001100110011010,
    22'b0000000100111101011100,
    22'b0000000001010001111011,
    22'b1111111110011001100110,
    22'b1111111101100110011010,
    22'b1111111101111010111000,
    22'b1111111111000010100100,
    22'b0000000000101000111101,
    22'b0000000011101011100001,
    22'b0000000110001111010111,
    22'b0000001000111101011100,
    22'b0000001011101011100001,
    22'b0000001101111010111000,
    22'b0000010000011110101110,
    22'b0000010010011001100110,
    22'b0000010011000010100100,
    22'b0000010010001111010111,
    22'b0000010000000000000000,
    22'b0000001101110000101001,
    22'b0000001011100001010010,
    22'b0000001001010001111011,
    22'b0000000111000010100100,
    22'b0000000100000000000000,
    22'b0000000010001111010111,
    22'b0000000000111101011100,
    22'b0000000000011110101110,
    22'b0000000000011110101110,
    22'b0000000001000111101100,
    22'b0000000001111010111000,
    22'b0000000010111000010100,
    22'b0000000011110101110001,
    22'b0000000101010001111011,
    22'b0000000110000101001000,
    22'b0000000110111000010100,
    22'b0000000111101011100001,
    22'b0000001000010100011111,
    22'b0000001000011110101110,
    22'b0000000111110101110001,
    22'b1111111110101110000101,
    22'b1111111010011001100110,
    22'b1111111001110000101001,
    22'b1111111000101000111101,
    22'b1111111001010001111011,
    22'b1111111100010100011111,
    22'b1111111111100001010010,
    22'b0000000010100011110110,
    22'b0000000101100110011010,
    22'b0000001001100110011010,
    22'b0000001100110011001101,
    22'b0000010000000000000000,
    22'b0000010011000010100100,
    22'b0000010101011100001010,
    22'b0000011000000000000000,
    22'b0000011001100110011010,
    22'b0000011010111000010100,
    22'b0000011100001010001111,
    22'b0000011101110000101001,
    22'b0000011111010111000011,
    22'b0000100001000111101100,
    22'b0000100010111000010100,
    22'b0000100100111101011100,
    22'b0000100110100011110110,
    22'b0000101000000000000000,
    22'b0000101001011100001010,
    22'b0000101011001100110011,
    22'b0000101101010001111011,
    22'b0000101111000010100100,
    22'b0000110000110011001101,
    22'b0000110011001100110011,
    22'b0000110101000111101100,
    22'b0000110101111010111000,
    22'b0000110110011001100110,
    22'b0000110110100011110110,
    22'b0000110110100011110110,
    22'b0000110110001111010111,
    22'b0000110101100110011010,
    22'b0000110100110011001101,
    22'b0000110011110101110001,
    22'b0000110011010111000011,
    22'b0000110010101110000101,
    22'b0000110010000101001000,
    22'b0000110001010001111011,
    22'b0000110000110011001101,
    22'b0000110000101000111101,
    22'b0000110000101000111101,
    22'b0000110000110011001101,
    22'b0000110000111101011100,
    22'b0000110000110011001101,
    22'b0000110000011110101110,
    22'b0000110000000000000000,
    22'b0000101111010111000011,
    22'b0000101111000010100100,
    22'b0000101110101110000101,
    22'b0000101110011001100110,
    22'b0000101101111010111000,
    22'b0000101101110000101001,
    22'b0000101101110000101001,
    22'b0000101101111010111000,
    22'b0000101101111010111000,
    22'b0000101110000101001000,
    22'b0000101110000101001000,
    22'b0000101110000101001000,
    22'b0000101101111010111000,
    22'b0000101101111010111000,
    22'b0000101101100110011010,
    22'b0000101100111101011100,
    22'b0000101100010100011111,
    22'b0000101011001100110011,
    22'b0000101010101110000101,
    22'b0000101010011001100110,
    22'b0000101010000101001000,
    22'b0000101001011100001010,
    22'b0000101000111101011100,
    22'b0000101000001010001111,
    22'b0000100111100001010010,
    22'b0000100110101110000101,
    22'b0000100110001111010111,
    22'b0000100101100110011010,
    22'b0000100100101000111101,
    22'b0000100101010001111011,
    22'b0000100101111010111000,
    22'b0000100110001111010111,
    22'b0000100110101110000101,
    22'b0000100110101110000101,
    22'b0000100110101110000101,
    22'b0000100110100011110110,
    22'b0000100110000101001000,
    22'b0000100101110000101001,
    22'b0000100101010001111011,
    22'b0000100100011110101110,
    22'b0000100011001100110011,
    22'b0000100010011001100110,
    22'b0000100001011100001010,
    22'b0000100000101000111101,
    22'b0000011111101011100001,
    22'b0000011110111000010100,
    22'b0000011110001111010111,
    22'b0000011101100110011010,
    22'b0000011100111101011100,
    22'b0000011100011110101110,
    22'b0000011011110101110001,
    22'b0000011011001100110011,
    22'b0000011010101110000101,
    22'b0000011010001111010111,
    22'b0000011001111010111000,
    22'b0000011001100110011010,
    22'b0000011001011100001010,
    22'b0000011001011100001010,
    22'b0000011001011100001010,
    22'b0000011001100110011010,
    22'b0000011010000101001000,
    22'b0000011010100011110110,
    22'b0000011011000010100100,
    22'b0000011011110101110001,
    22'b0000011100010100011111,
    22'b0000011101010001111011,
    22'b0000011111100001010010,
    22'b0000100001110000101001,
    22'b0000100001100110011010,
    22'b0000100000101000111101,
    22'b0000011100010100011111,
    22'b0000011011010111000011,
    22'b0000011010100011110110,
    22'b0000011010000101001000,
    22'b0000011010000101001000,
    22'b0000011010100011110110,
    22'b0000011011001100110011,
    22'b0000011100001010001111,
    22'b0000011101111010111000,
    22'b0000011110111000010100,
    22'b0000011111110101110001,
    22'b0000100000111101011100,
    22'b0000100001100110011010,
    22'b0000100010000101001000,
    22'b0000100010011001100110,
    22'b0000100010111000010100,
    22'b0000100010111000010100,
    22'b0000100010100011110110,
    22'b0000100010000101001000,
    22'b0000100001010001111011,
    22'b0000100000011110101110,
    22'b0000011111101011100001,
    22'b0000011110111000010100,
    22'b0000011110000101001000,
    22'b0000011101100110011010,
    22'b0000011101000111101100,
    22'b0000011100110011001101,
    22'b0000011100011110101110,
    22'b0000011100010100011111,
    22'b0000011100000000000000,
    22'b0000011011110101110001,
    22'b0000011011110101110001,
    22'b0000011100000000000000,
    22'b0000011101010001111011,
    22'b0000011101000111101100,
    22'b0000011100101000111101,
    22'b0000011100010100011111,
    22'b0000011100010100011111,
    22'b0000011100001010001111,
    22'b0000011100001010001111,
    22'b0000011100001010001111,
    22'b0000011100010100011111,
    22'b0000011100111101011100,
    22'b0000011101110000101001,
    22'b0000011110111000010100,
    22'b0000011111001100110011,
    22'b0000011111010111000011,
    22'b0000011111101011100001,
    22'b0000011111100001010010,
    22'b0000011111010111000011,
    22'b0000011111001100110011,
    22'b0000011110111000010100,
    22'b0000011110011001100110,
    22'b0000011101111010111000,
    22'b0000011100111101011100,
    22'b0000011011101011100001,
    22'b0000011010100011110110,
    22'b0000011001010001111011,
    22'b0000010111100001010010,
    22'b0000010110000101001000,
    22'b0000010100110011001101,
    22'b0000010011110101110001,
    22'b0000010011010111000011,
    22'b0000010011101011100001,
    22'b0000010110001111010111,
    22'b0000010110011001100110,
    22'b0000010110001111010111,
    22'b0000010101111010111000,
    22'b0000010101010001111011,
    22'b0000010100101000111101,
    22'b0000010100000000000000,
    22'b0000010011001100110011,
    22'b0000010010001111010111,
    22'b0000010001100110011010,
    22'b0000010000110011001101,
    22'b0000010000000000000000,
    22'b0000001111000010100100,
    22'b0000001110100011110110,
    22'b0000001101111010111000,
    22'b0000001101010001111011,
    22'b0000001100110011001101,
    22'b0000001100011110101110,
    22'b0000001100001010001111,
    22'b0000001011101011100001,
    22'b0000001011001100110011,
    22'b0000001010111000010100,
    22'b0000001010100011110110,
    22'b0000001010011001100110,
    22'b0000001010001111010111,
    22'b0000001010000101001000,
    22'b0000001010001111010111,
    22'b0000001010100011110110,
    22'b0000001011010111000011,
    22'b0000001100010100011111,
    22'b0000001101111010111000,
    22'b0000010100011110101110,
    22'b0000010110011001100110,
    22'b0000011000001010001111,
    22'b0000011000111101011100,
    22'b0000011001011100001010,
    22'b0000011001010001111011,
    22'b0000011000110011001101,
    22'b0000011000001010001111,
    22'b0000010111100001010010,
    22'b0000010110100011110110,
    22'b0000010101111010111000,
    22'b0000010101010001111011,
    22'b0000010100010100011111,
    22'b0000010010101110000101,
    22'b0000010001010001111011,
    22'b0000001111110101110001,
    22'b0000001110000101001000,
    22'b0000001100101000111101,
    22'b0000001011010111000011,
    22'b0000001010000101001000,
    22'b0000001000001010001111,
    22'b0000000110100011110110,
    22'b0000000100111101011100,
    22'b0000000011001100110011,
    22'b0000000001000111101100,
    22'b1111111111101011100001,
    22'b1111111110001111010111,
    22'b1111111100011110101110,
    22'b1111111011100001010010,
    22'b1111111010100011110110,
    22'b1111111001110000101001,
    22'b1111111000110011001101,
    22'b1111111000101000111101,
    22'b1111111000101000111101,
    22'b1111111000101000111101,
    22'b1111111000101000111101,
    22'b1111111000110011001101,
    22'b1111111000110011001101,
    22'b1111111000110011001101,
    22'b1111111000110011001101,
    22'b1111111000101000111101,
    22'b1111111000011110101110,
    22'b1111111000010100011111,
    22'b1111111000000000000000,
    22'b1111110111101011100001,
    22'b1111110111001100110011,
    22'b1111110110111000010100,
    22'b1111110110100011110110,
    22'b1111110110100011110110,
    22'b1111110110111000010100,
    22'b1111110111100001010010,
    22'b1111111000011110101110,
    22'b1111111001111010111000,
    22'b1111111011000010100100,
    22'b1111111100010100011111,
    22'b1111111110011001100110,
    22'b1111111111101011100001,
    22'b0000000000110011001101,
    22'b0000000001011100001010,
    22'b0000000001111010111000,
    22'b0000000001111010111000,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001000111101100,
    22'b0000000000110011001101,
    22'b0000000000101000111101,
    22'b0000000000011110101110,
    22'b0000000000110011001101,
    22'b0000000001010001111011,
    22'b0000000001111010111000,
    22'b0000000010101110000101,
    22'b0000000100000000000000,
    22'b0000000101000111101100,
    22'b0000000101111010111000,
    22'b0000000111001100110011,
    22'b0000001000001010001111,
    22'b0000001001000111101100,
    22'b0000001010000101001000,
    22'b0000001011100001010010,
    22'b0000001100010100011111,
    22'b0000001100111101011100,
    22'b0000001101110000101001,
    22'b0000001110011001100110,
    22'b0000001110111000010100,
    22'b0000001111000010100100,
    22'b0000001110101110000101,
    22'b0000001101110000101001,
    22'b0000001100110011001101,
    22'b0000001011110101110001,
    22'b0000001010101110000101,
    22'b0000001001111010111000,
    22'b0000000110000101001000,
    22'b0000000100111101011100,
    22'b0000000100010100011111,
    22'b0000000011110101110001,
    22'b0000000011100001010010,
    22'b0000000011010111000011,
    22'b0000000011001100110011,
    22'b0000000011001100110011,
    22'b0000000011001100110011,
    22'b0000000011001100110011,
    22'b0000000011001100110011,
    22'b0000000011000010100100,
    22'b0000000010111000010100,
    22'b0000000010011001100110,
    22'b0000000001110000101001,
    22'b0000000000110011001101,
    22'b1111111111101011100001,
    22'b1111111110101110000101,
    22'b1111111110000101001000,
    22'b1111111110000101001000,
    22'b1111111110001111010111,
    22'b1111111110100011110110,
    22'b1111111111000010100100,
    22'b1111111111101011100001,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111110011001100110,
    22'b1111111101111010111000,
    22'b1111111101010001111011,
    22'b1111111110001111010111,
    22'b1111111111010111000011,
    22'b0000000000011110101110,
    22'b0000000010001111010111,
    22'b0000000011101011100001,
    22'b0000000101000111101100,
    22'b0000000110011001100110,
    22'b0000001000000000000000,
    22'b0000001001010001111011,
    22'b0000001010100011110110,
    22'b0000001011101011100001,
    22'b0000001100011110101110,
    22'b0000001100111101011100,
    22'b0000001101111010111000,
    22'b0000001110111000010100,
    22'b0000001111001100110011,
    22'b0000001111001100110011,
    22'b0000001111101011100001,
    22'b0000001111001100110011,
    22'b0000001110101110000101,
    22'b0000001110011001100110,
    22'b0000001110100011110110,
    22'b0000001110111000010100,
    22'b0000001110111000010100,
    22'b0000001110000101001000,
    22'b0000001100110011001101,
    22'b0000001011110101110001,
    22'b0000001100011110101110,
    22'b0000001101011100001010,
    22'b0000010001011100001010,
    22'b0000010001000111101100,
    22'b0000010000110011001101,
    22'b0000010000010100011111,
    22'b0000001111010111000011,
    22'b0000001110011001100110,
    22'b0000001101011100001010,
    22'b0000001100001010001111,
    22'b0000001100101000111101,
    22'b0000001100111101011100,
    22'b0000001100110011001101,
    22'b0000001100110011001101,
    22'b0000001100101000111101,
    22'b0000001100101000111101,
    22'b0000001101010001111011,
    22'b0000001101111010111000,
    22'b0000001110001111010111,
    22'b0000001110000101001000,
    22'b0000001101111010111000,
    22'b0000001101000111101100,
    22'b0000001100010100011111,
    22'b0000001010111000010100,
    22'b0000001000111101011100,
    22'b0000000111000010100100,
    22'b0000000100111101011100,
    22'b0000000100001010001111,
    22'b0000000100110011001101,
    22'b0000000110011001100110,
    22'b0000001000101000111101,
    22'b0000001010001111010111,
    22'b0000001010000101001000,
    22'b0000000111110101110001,
    22'b0000000100111101011100,
    22'b0000000010101110000101,
    22'b0000000001110000101001,
    22'b0000000011000010100100,
    22'b0000000100010100011111,
    22'b0000000100011110101110,
    22'b0000000011101011100001,
    22'b0000000011110101110001,
    22'b0000000011001100110011,
    22'b0000000011101011100001,
    22'b0000000011110101110001,
    22'b0000000100001010001111,
    22'b0000000011101011100001,
    22'b0000000010101110000101,
    22'b0000000011001100110011,
    22'b0000000010101110000101,
    22'b0000000011101011100001,
    22'b0000000011100001010010,
    22'b0000000011100001010010,
    22'b0000000100101000111101,
    22'b0000000100111101011100,
    22'b0000000110001111010111,
    22'b0000000101110000101001,
    22'b0000000101000111101100,
    22'b0000000100011110101110,
    22'b0000000100101000111101,
    22'b0000000101100110011010,
    22'b0000000101110000101001,
    22'b0000000101011100001010,
    22'b0000000001000111101100,
    22'b0000000000110011001101,
    22'b0000000000001010001111,
    22'b1111111111101011100001,
    22'b1111111111010111000011,
    22'b1111111111010111000011,
    22'b1111111111001100110011,
    22'b1111111111001100110011,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111010111000011,
    22'b1111111110111000010100,
    22'b1111111110011001100110,
    22'b1111111110000101001000,
    22'b1111111101110000101001,
    22'b1111111101110000101001,
    22'b1111111110000101001000,
    22'b1111111110101110000101,
    22'b1111111111100001010010,
    22'b0000000000111101011100,
    22'b0000000010000101001000,
    22'b0000000011000010100100,
    22'b0000000011110101110001,
    22'b0000000100011110101110,
    22'b0000000100110011001101,
    22'b0000000100111101011100,
    22'b0000000101000111101100,
    22'b0000000100111101011100,
    22'b0000000100110011001101,
    22'b0000000100001010001111,
    22'b0000000011000010100100,
    22'b0000000001000111101100,
    22'b1111111111010111000011,
    22'b1111111101011100001010,
    22'b1111111011010111000011,
    22'b1111111000111101011100,
    22'b1111101110100011110110,
    22'b1111101100111101011100,
    22'b1111101011000010100100,
    22'b1111101000101000111101,
    22'b1111100111001100110011,
    22'b1111100111100001010010,
    22'b1111101000011110101110,
    22'b1111101010101110000101,
    22'b1111101100011110101110,
    22'b1111101101100110011010,
    22'b1111101110100011110110,
    22'b1111101111110101110001,
    22'b1111110001000111101100,
    22'b1111110010111000010100,
    22'b1111110100101000111101,
    22'b1111110111000010100100,
    22'b1111111000010100011111,
    22'b1111111001000111101100,
    22'b1111111001100110011010,
    22'b1111111001111010111000,
    22'b1111111010000101001000,
    22'b1111111001111010111000,
    22'b1111111001100110011010,
    22'b1111111000101000111101,
    22'b1111110111100001010010,
    22'b1111110110001111010111,
    22'b1111110100110011001101,
    22'b1111110010100011110110,
    22'b1111110000110011001101,
    22'b1111101110111000010100,
    22'b1111101100110011001101,
    22'b1111101001111010111000,
    22'b1111100111110101110001,
    22'b1111100110000101001000,
    22'b1111100100010100011111,
    22'b1111100010001111010111,
    22'b1111100000110011001101,
    22'b1111011100011110101110,
    22'b1111011101010001111011,
    22'b1111100000000000000000,
    22'b1111100011010111000011,
    22'b1111100111100001010010,
    22'b1111101011110101110001,
    22'b1111110000110011001101,
    22'b1111110011110101110001,
    22'b1111110110000101001000,
    22'b1111110111100001010010,
    22'b1111111000110011001101,
    22'b1111111001000111101100,
    22'b1111111001011100001010,
    22'b1111111001011100001010,
    22'b1111111001000111101100,
    22'b1111111000011110101110,
    22'b1111110111101011100001,
    22'b1111110110101110000101,
    22'b1111110101010001111011,
    22'b1111110100001010001111,
    22'b1111110011001100110011,
    22'b1111110010100011110110,
    22'b1111110010000101001000,
    22'b1111110001110000101001,
    22'b1111110001100110011010,
    22'b1111110001011100001010,
    22'b1111110001000111101100,
    22'b1111110000110011001101,
    22'b1111110000011110101110,
    22'b1111110000000000000000,
    22'b1111101111001100110011,
    22'b1111101110011001100110,
    22'b1111101101100110011010,
    22'b1111101100110011001101,
    22'b1111101100000000000000,
    22'b1111101010111000010100,
    22'b1111101010001111010111,
    22'b1111101001110000101001,
    22'b1111101010000101001000,
    22'b1111110010000101001000,
    22'b1111110011101011100001,
    22'b1111110100111101011100,
    22'b1111110110011001100110,
    22'b1111110111001100110011,
    22'b1111110111110101110001,
    22'b1111111000010100011111,
    22'b1111111000101000111101,
    22'b1111111000101000111101,
    22'b1111111000011110101110,
    22'b1111111000001010001111,
    22'b1111110111100001010010,
    22'b1111110111001100110011,
    22'b1111110110101110000101,
    22'b1111110110011001100110,
    22'b1111110110000101001000,
    22'b1111110101110000101001,
    22'b1111110101010001111011,
    22'b1111110100011110101110,
    22'b1111110011101011100001,
    22'b1111110010111000010100,
    22'b1111110001110000101001,
    22'b1111110000001010001111,
    22'b1111101110111000010100,
    22'b1111101101110000101001,
    22'b1111101100011110101110,
    22'b1111101010111000010100,
    22'b1111101001110000101001,
    22'b1111101000110011001101,
    22'b1111100111101011100001,
    22'b1111100110000101001000,
    22'b1111100100111101011100,
    22'b1111100011101011100001,
    22'b1111100010100011110110,
    22'b1111100000101000111101,
    22'b1111011111001100110011,
    22'b1111011110001111010111,
    22'b1111011101010001111011,
    22'b1111011100110011001101,
    22'b1111011100011110101110,
    22'b1111011100010100011111,
    22'b1111011100001010001111,
    22'b1111011101000111101100,
    22'b1111011101111010111000,
    22'b1111011111001100110011,
    22'b1111100000010100011111,
    22'b1111100001011100001010,
    22'b1111100010100011110110,
    22'b1111100100010100011111,
    22'b1111100101110000101001,
    22'b1111100111010111000011,
    22'b1111101000110011001101,
    22'b1111101010101110000101,
    22'b1111101011110101110001,
    22'b1111101100110011001101,
    22'b1111101101100110011010,
    22'b1111101110001111010111,
    22'b1111101110100011110110,
    22'b1111101110111000010100,
    22'b1111101111000010100100,
    22'b1111101111001100110011,
    22'b1111101111001100110011,
    22'b1111101111001100110011,
    22'b1111101111000010100100,
    22'b1111101110111000010100,
    22'b1111101110101110000101,
    22'b1111101110011001100110,
    22'b1111101110001111010111,
    22'b1111101101111010111000,
    22'b1111101101100110011010,
    22'b1111101101011100001010,
    22'b1111101101000111101100,
    22'b1111101100101000111101,
    22'b1111101100011110101110,
    22'b1111101100010100011111,
    22'b1111101100001010001111,
    22'b1111101100001010001111,
    22'b1111101100010100011111,
    22'b1111101100101000111101,
    22'b1111101101000111101100,
    22'b1111101110000101001000,
    22'b1111101110111000010100,
    22'b1111110000000000000000,
    22'b1111110001000111101100,
    22'b1111110010000101001000,
    22'b1111110011000010100100,
    22'b1111110011010111000011,
    22'b1111110011110101110001,
    22'b1111110100011110101110,
    22'b1111110101100110011010,
    22'b1111110110100011110110,
    22'b1111110111110101110001,
    22'b1111111001000111101100,
    22'b1111111001010001111011,
    22'b1111111001100110011010,
    22'b1111111010111000010100,
    22'b1111111100110011001101,
    22'b1111111101010001111011,
    22'b1111111011010111000011,
    22'b1111111010101110000101,
    22'b1111111001110000101001,
    22'b1111111000111101011100,
    22'b1111111000011110101110,
    22'b1111111000011110101110,
    22'b1111110111000010100100,
    22'b1111110101110000101001,
    22'b1111110100010100011111,
    22'b1111110011010111000011,
    22'b1111110010011001100110,
    22'b1111110001100110011010,
    22'b1111110001010001111011,
    22'b1111110000111101011100,
    22'b1111110000111101011100,
    22'b1111110001000111101100,
    22'b1111110001011100001010,
    22'b1111110010000101001000,
    22'b1111110011100001010010,
    22'b1111111000011110101110,
    22'b1111111010011001100110,
    22'b1111111001111010111000,
    22'b1111111000111101011100,
    22'b1111111000010100011111,
    22'b1111110111110101110001,
    22'b1111111000001010001111,
    22'b1111111000110011001101,
    22'b1111111001000111101100,
    22'b1111111001000111101100,
    22'b1111111000110011001101,
    22'b1111111000101000111101,
    22'b1111111000011110101110,
    22'b1111111000101000111101,
    22'b1111111001000111101100,
    22'b1111111001100110011010,
    22'b1111111010001111010111,
    22'b1111111010111000010100,
    22'b1111111011010111000011,
    22'b1111111011000010100100,
    22'b1111111010011001100110,
    22'b1111111001000111101100,
    22'b1111110111010111000011,
    22'b1111110100111101011100,
    22'b1111110011010111000011,
    22'b1111110001111010111000,
    22'b1111110000110011001101,
    22'b1111101111001100110011,
    22'b1111101110001111010111,
    22'b1111101101011100001010,
    22'b1111101101010001111011,
    22'b1111101101111010111000,
    22'b1111101111000010100100,
    22'b1111110000110011001101,
    22'b1111110010111000010100,
    22'b1111110101010001111011,
    22'b1111110111100001010010,
    22'b1111111000000000000000,
    22'b1111111000110011001101,
    22'b1111111001010001111011,
    22'b1111111001011100001010,
    22'b1111111001110000101001,
    22'b1111111001110000101001,
    22'b1111111010000101001000,
    22'b1111111001111010111000,
    22'b1111111001011100001010,
    22'b1111111001110000101001,
    22'b1111111000110011001101,
    22'b1111111000101000111101,
    22'b1111111001110000101001,
    22'b1111111010011001100110,
    22'b1111111010011001100110,
    22'b1111111010100011110110,
    22'b1111111011000010100100,
    22'b1111111011100001010010,
    22'b1111111011110101110001,
    22'b1111111100001010001111,
    22'b1111111100010100011111,
    22'b1111111100000000000000,
    22'b1111111011100001010010,
    22'b1111111011001100110011,
    22'b1111111011010111000011,
    22'b1111111011010111000011,
    22'b1111111011101011100001,
    22'b1111111100000000000000,
    22'b1111111100111101011100,
    22'b1111111110100011110110,
    22'b0000000000000000000000,
    22'b0000000000110011001101,
    22'b0000000001110000101001,
    22'b0000000011001100110011,
    22'b0000000100101000111101,
    22'b0000000101011100001010,
    22'b0000000101111010111000,
    22'b0000000101100110011010,
    22'b0000000101000111101100,
    22'b0000000100011110101110,
    22'b0000000011101011100001,
    22'b0000000011000010100100,
    22'b0000000010000101001000,
    22'b0000000001011100001010,
    22'b0000000000101000111101,
    22'b1111111111110101110001,
    22'b1111111111100001010010,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111101011100001,
    22'b1111111111110101110001,
    22'b0000000001111010111000,
    22'b0000000010011001100110,
    22'b0000000011000010100100,
    22'b0000000100001010001111,
    22'b0000000101100110011010,
    22'b0000000111010111000011,
    22'b0000001000111101011100,
    22'b0000001010100011110110,
    22'b0000001100011110101110,
    22'b0000001101111010111000,
    22'b0000001111001100110011,
    22'b0000010000011110101110,
    22'b0000010001110000101001,
    22'b0000010010100011110110,
    22'b0000010011001100110011,
    22'b0000010011110101110001,
    22'b0000010100001010001111,
    22'b0000010100001010001111,
    22'b0000010101000111101100,
    22'b0000010101110000101001,
    22'b0000010110111000010100,
    22'b0000011000010100011111,
    22'b0000011001011100001010,
    22'b0000011010001111010111,
    22'b0000011011001100110011,
    22'b0000011100000000000000,
    22'b0000011100111101011100,
    22'b0000011101010001111011,
    22'b0000011101110000101001,
    22'b0000011110000101001000,
    22'b0000011110011001100110,
    22'b0000011111101011100001,
    22'b0000100000101000111101,
    22'b0000100001100110011010,
    22'b0000100010011001100110,
    22'b0000100010101110000101,
    22'b0000100010111000010100,
    22'b0000100010100011110110,
    22'b0000100010101110000101,
    22'b0000100010111000010100,
    22'b0000100011100001010010,
    22'b0000100100101000111101,
    22'b0000100101011100001010,
    22'b0000100101011100001010,
    22'b0000100100111101011100,
    22'b0000100100011110101110,
    22'b0000100100001010001111,
    22'b0000100100001010001111,
    22'b0000100100010100011111,
    22'b0000100100011110101110,
    22'b0000100100111101011100,
    22'b0000100100111101011100,
    22'b0000100101000111101100,
    22'b0000100100101000111101,
    22'b0000100100001010001111,
    22'b0000100011010111000011,
    22'b0000100010100011110110,
    22'b0000100001010001111011,
    22'b0000011110111000010100,
    22'b0000011100111101011100,
    22'b0000011011001100110011,
    22'b0000011001111010111000,
    22'b0000011000110011001101,
    22'b0000011000010100011111,
    22'b0000010111101011100001,
    22'b0000010111001100110011,
    22'b0000010110111000010100,
    22'b0000010110001111010111,
    22'b0000010101100110011010,
    22'b0000010101011100001010,
    22'b0000010101000111101100,
    22'b0000010101000111101100,
    22'b0000010101010001111011,
    22'b0000010101011100001010,
    22'b0000010101011100001010,
    22'b0000010101011100001010,
    22'b0000010101010001111011,
    22'b0000010100111101011100,
    22'b0000010100101000111101,
    22'b0000010100001010001111,
    22'b0000010011100001010010,
    22'b0000010011000010100100,
    22'b0000010010001111010111,
    22'b0000010001010001111011,
    22'b0000010000000000000000,
    22'b0000001100111101011100,
    22'b0000001100011110101110,
    22'b0000001100001010001111,
    22'b0000001011101011100001,
    22'b0000001011100001010010,
    22'b0000001011010111000011,
    22'b0000001011000010100100,
    22'b0000001010001111010111,
    22'b0000001000111101011100,
    22'b0000000111010111000011,
    22'b0000000100101000111101,
    22'b0000000010011001100110,
    22'b1111111111010111000011,
    22'b1111111100111101011100,
    22'b1111111100011110101110,
    22'b1111111010101110000101,
    22'b1111111010001111010111,
    22'b1111111010100011110110,
    22'b1111111010100011110110,
    22'b1111111010111000010100,
    22'b1111111100000000000000,
    22'b1111111100010100011111,
    22'b1111111100011110101110,
    22'b1111111100011110101110,
    22'b1111111100000000000000,
    22'b1111111010101110000101,
    22'b1111111001100110011010,
    22'b1111110111010111000011,
    22'b1111110100011110101110,
    22'b1111110010000101001000,
    22'b1111101111001100110011,
    22'b1111101100011110101110,
    22'b1111100111010111000011,
    22'b1111100100101000111101,
    22'b1111100000111101011100,
    22'b1111011101011100001010,
    22'b1111011011000010100100,
    22'b1111011010011001100110,
    22'b1111011010011001100110,
    22'b1111011001100110011010,
    22'b1111011001000111101100,
    22'b1111011000110011001101,
    22'b1111011001000111101100,
    22'b1111011000110011001101,
    22'b1111011000101000111101,
    22'b1111010111101011100001,
    22'b1111010110100011110110,
    22'b1111010111000010100100,
    22'b1111010111001100110011,
    22'b1111010111100001010010,
    22'b1111010110111000010100,
    22'b1111010111101011100001,
    22'b1111011001000111101100,
    22'b1111011010011001100110,
    22'b1111011011001100110011,
    22'b1111011100110011001101,
    22'b1111011110100011110110,
    22'b1111011111110101110001,
    22'b1111100000101000111101,
    22'b1111100001110000101001,
    22'b1111100010011001100110,
    22'b1111100011001100110011,
    22'b1111100100101000111101,
    22'b1111100101100110011010,
    22'b1111100110011001100110,
    22'b1111100110001111010111,
    22'b1111100110111000010100,
    22'b1111100110011001100110,
    22'b1111101000000000000000,
    22'b1111100110111000010100,
    22'b1111100110000101001000,
    22'b1111100001010001111011,
    22'b1111011010000101001000,
    22'b1111010100001010001111,
    22'b1111001110001111010111,
    22'b1111001001111010111000,
    22'b1111000110011001100110,
    22'b1111000100110011001101,
    22'b1111000100110011001101,
    22'b1111000110000101001000,
    22'b1111001001011100001010,
    22'b1111001100011110101110,
    22'b1111001111101011100001,
    22'b1111010011000010100100,
    22'b1111010111101011100001,
    22'b1111011010100011110110,
    22'b1111011100101000111101,
    22'b1111011111000010100100,
    22'b1111100000101000111101,
    22'b1111100001111010111000,
    22'b1111100011010111000011,
    22'b1111100101100110011010,
    22'b1111100111101011100001,
    22'b1111101001100110011010,
    22'b1111101111100001010010,
    22'b1111101111100001010010,
    22'b1111101111010111000011,
    22'b1111101110001111010111,
    22'b1111101101000111101100,
    22'b1111101100000000000000,
    22'b1111101010011001100110,
    22'b1111101000000000000000,
    22'b1111100110001111010111,
    22'b1111100100011110101110,
    22'b1111100010101110000101,
    22'b1111100001110000101001,
    22'b1111100000101000111101,
    22'b1111011111101011100001,
    22'b1111011111100001010010,
    22'b1111011111100001010010,
    22'b1111100000011110101110,
    22'b1111100010000101001000,
    22'b1111100100110011001101,
    22'b1111100111001100110011,
    22'b1111101010101110000101,
    22'b1111101110101110000101,
    22'b1111110001000111101100,
    22'b1111110011110101110001,
    22'b1111110101110000101001,
    22'b1111111000000000000000,
    22'b1111111001010001111011,
    22'b1111111010100011110110,
    22'b1111111011100001010010,
    22'b1111111101000111101100,
    22'b0000000011110101110001,
    22'b0000000101100110011010,
    22'b0000000111100001010010,
    22'b0000001000101000111101,
    22'b0000001001100110011010,
    22'b0000001010000101001000,
    22'b0000001001111010111000,
    22'b0000001001011100001010,
    22'b0000001000011110101110,
    22'b0000000110101110000101,
    22'b0000000101000111101100,
    22'b0000000011010111000011,
    22'b0000000001010001111011,
    22'b1111111110011001100110,
    22'b1111111100011110101110,
    22'b1111111010111000010100,
    22'b1111111001100110011010,
    22'b1111111000010100011111,
    22'b1111110111110101110001,
    22'b1111110111100001010010,
    22'b1111110111001100110011,
    22'b1111110111000010100100,
    22'b1111110110101110000101,
    22'b1111110110101110000101,
    22'b1111110110111000010100,
    22'b1111110110111000010100,
    22'b1111110111000010100100,
    22'b1111110111010111000011,
    22'b1111111000110011001101,
    22'b1111111001110000101001,
    22'b1111111010111000010100,
    22'b1111111100000000000000,
    22'b1111111101011100001010,
    22'b1111111110011001100110,
    22'b1111111111100001010010,
    22'b0000000101010001111011,
    22'b0000000110001111010111,
    22'b0000000110011001100110,
    22'b0000000110001111010111,
    22'b0000000110011001100110,
    22'b0000000110011001100110,
    22'b0000000110000101001000,
    22'b0000000110000101001000,
    22'b0000000110001111010111,
    22'b0000000110011001100110,
    22'b0000000110100011110110,
    22'b0000000111000010100100,
    22'b0000000111100001010010,
    22'b0000000111110101110001,
    22'b0000001000010100011111,
    22'b0000001001010001111011,
    22'b0000001001111010111000,
    22'b0000001010101110000101,
    22'b0000001011101011100001,
    22'b0000001100110011001101,
    22'b0000001101110000101001,
    22'b0000001110111000010100,
    22'b0000010000011110101110,
    22'b0000010010000101001000,
    22'b0000010011101011100001,
    22'b0000010101011100001010,
    22'b0000010111110101110001,
    22'b0000011001100110011010,
    22'b0000011011001100110011,
    22'b0000011100101000111101,
    22'b0000011110011001100110,
    22'b0000011111101011100001,
    22'b0000100000011110101110,
    22'b0000100001010001111011,
    22'b0000100001110000101001,
    22'b0000100001100110011010,
    22'b0000100000110011001101,
    22'b0000011111101011100001,
    22'b0000011101010001111011,
    22'b0000011010111000010100,
    22'b0000011000010100011111,
    22'b0000010110000101001000,
    22'b0000001101011100001010,
    22'b0000001100011110101110,
    22'b0000001100001010001111,
    22'b0000001100000000000000,
    22'b0000001011100001010010,
    22'b0000001010000101001000,
    22'b0000001001010001111011,
    22'b0000001000010100011111,
    22'b0000001000000000000000,
    22'b0000000111001100110011,
    22'b0000000101010001111011,
    22'b0000000100010100011111,
    22'b0000000011000010100100,
    22'b0000000010001111010111,
    22'b0000000001111010111000,
    22'b0000000000110011001101,
    22'b1111111110100011110110,
    22'b1111111100111101011100,
    22'b1111111100000000000000,
    22'b1111111001000111101100,
    22'b1111110110100011110110,
    22'b1111110100110011001101,
    22'b1111110001010001111011,
    22'b1111101110000101001000,
    22'b1111101011000010100100,
    22'b1111101000001010001111,
    22'b1111100011101011100001,
    22'b1111011111100001010010,
    22'b1111011010101110000101,
    22'b1111010101000111101100,
    22'b1111001101110000101001,
    22'b1111001001110000101001,
    22'b1111000101110000101001,
    22'b1111000000011110101110,
    22'b1110111100111101011100,
    22'b1110111010000101001000,
    22'b1110110111101011100001,
    22'b1110110110100011110110,
    22'b1110111000010100011111,
    22'b1111001010100011110110,
    22'b1111010001010001111011,
    22'b1111010101100110011010,
    22'b1111011001100110011010,
    22'b1111011100101000111101,
    22'b1111011111110101110001,
    22'b1111100001100110011010,
    22'b1111100011010111000011,
    22'b1111100101010001111011,
    22'b1111100110100011110110,
    22'b1111100111110101110001,
    22'b1111101000110011001101,
    22'b1111101010011001100110,
    22'b1111101011100001010010,
    22'b1111101100110011001101,
    22'b1111101110011001100110,
    22'b1111101111010111000011,
    22'b1111110000000000000000,
    22'b1111110000001010001111,
    22'b1111110000000000000000,
    22'b1111101111010111000011,
    22'b1111101101111010111000,
    22'b1111101100001010001111,
    22'b1111101001000111101100,
    22'b1111100111000010100100,
    22'b1111100100011110101110,
    22'b1111100001100110011010,
    22'b1111011111101011100001,
    22'b1111011110001111010111,
    22'b1111011101100110011010,
    22'b1111011101000111101100,
    22'b1111011100000000000000,
    22'b1111011010001111010111,
    22'b1111011001100110011010,
    22'b1111010101000111101100,
    22'b1111011001000111101100,
    22'b1111011110100011110110,
    22'b1111100100001010001111,
    22'b1111101000111101011100,
    22'b1111101110000101001000,
    22'b1111110011001100110011,
    22'b1111111001000111101100,
    22'b1111111100010100011111,
    22'b1111111110000101001000,
    22'b1111111110111000010100,
    22'b1111111111000010100100,
    22'b1111111110101110000101,
    22'b1111111110100011110110,
    22'b1111111110101110000101,
    22'b1111111111000010100100,
    22'b1111111111001100110011,
    22'b1111111111010111000011,
    22'b1111111111101011100001,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111010111000011,
    22'b1111111110011001100110,
    22'b1111111100110011001101,
    22'b1111111011000010100100,
    22'b1111111001000111101100,
    22'b1111110111101011100001,
    22'b1111111000011110101110,
    22'b1111111011001100110011,
    22'b1111111101000111101100,
    22'b1111111101010001111011,
    22'b1111111100010100011111,
    22'b1111111010101110000101,
    22'b1111110111110101110001,
    22'b1111111001011100001010,
    22'b1111111100010100011111,
    22'b1111111111010111000011,
    22'b0000000000000000000000,
    22'b0000000000111101011100,
    22'b0000000001010001111011,
    22'b0000000001110000101001,
    22'b0000000011000010100100,
    22'b0000000011010111000011,
    22'b0000000100001010001111,
    22'b0000000011100001010010,
    22'b0000000011101011100001,
    22'b0000000101110000101001,
    22'b0000000100110011001101,
    22'b0000000100011110101110,
    22'b0000000101011100001010,
    22'b0000000100110011001101,
    22'b0000000100011110101110,
    22'b0000000101000111101100,
    22'b0000000000011110101110,
    22'b1111111000001010001111,
    22'b1111101101100110011010,
    22'b1111100101100110011010,
    22'b1111011010001111010111,
    22'b1111001001011100001010,
    22'b1111000010011001100110,
    22'b1110111011001100110011,
    22'b1110110100110011001101,
    22'b1110110011110101110001,
    22'b1110111001100110011010,
    22'b1111000000101000111101,
    22'b1111000111001100110011,
    22'b1111011000101000111101,
    22'b1111100100001010001111,
    22'b1111101101100110011010,
    22'b1111110110101110000101,
    22'b1111111011000010100100,
    22'b1111111010011001100110,
    22'b1111111010011001100110,
    22'b1111111011000010100100,
    22'b1111111100000000000000,
    22'b1111111101000111101100,
    22'b1111111110011001100110,
    22'b1111111111001100110011,
    22'b0000000000000000000000,
    22'b0000000000111101011100,
    22'b0000000001111010111000,
    22'b0000000011001100110011,
    22'b0000000100110011001101,
    22'b0000000111110101110001,
    22'b0000001010001111010111,
    22'b0000001100011110101110,
    22'b0000001110101110000101,
    22'b0000010000111101011100,
    22'b0000010010000101001000,
    22'b0000010011000010100100,
    22'b0000010011010111000011,
    22'b0000010010111000010100,
    22'b0000010001111010111000,
    22'b0000010000011110101110,
    22'b0000001110100011110110,
    22'b0000001101010001111011,
    22'b0000001100010100011111,
    22'b0000001011100001010010,
    22'b0000001010111000010100,
    22'b0000001010101110000101,
    22'b0000001010100011110110,
    22'b0000001010100011110110,
    22'b0000001100001010001111,
    22'b0000001100111101011100,
    22'b0000001101100110011010,
    22'b0000001101110000101001,
    22'b0000001101111010111000,
    22'b0000001101011100001010,
    22'b0000001100111101011100,
    22'b0000001100001010001111,
    22'b0000001011010111000011,
    22'b0000001011001100110011,
    22'b0000001100000000000000,
    22'b0000001101000111101100,
    22'b0000001110001111010111,
    22'b0000001111110101110001,
    22'b0000010000111101011100,
    22'b0000010010000101001000,
    22'b0000010011010111000011,
    22'b0000010101000111101100,
    22'b0000010110001111010111,
    22'b0000010111001100110011,
    22'b0000010111110101110001,
    22'b0000010111110101110001,
    22'b0000010110111000010100,
    22'b0000010101000111101100,
    22'b0000001110111000010100,
    22'b0000001010000101001000,
    22'b0000000111101011100001,
    22'b0000000101100110011010,
    22'b1111111110111000010100,
    22'b1111111100111101011100,
    22'b1111111101110000101001,
    22'b0000000100110011001101,
    22'b0000000110111000010100,
    22'b0000001000110011001101,
    22'b0000001010001111010111,
    22'b0000001011101011100001,
    22'b0000001100101000111101,
    22'b0000001101100110011010,
    22'b0000001110111000010100,
    22'b0000001101100110011010,
    22'b0000001101100110011010,
    22'b0000001111001100110011,
    22'b0000010000001010001111,
    22'b0000010000101000111101,
    22'b0000010010000101001000,
    22'b0000010011001100110011,
    22'b0000010101100110011010,
    22'b0000010111100001010010,
    22'b0000011000010100011111,
    22'b0000011000001010001111,
    22'b0000011000101000111101,
    22'b0000011000111101011100,
    22'b0000010111100001010010,
    22'b0000010010111000010100,
    22'b0000010010000101001000,
    22'b0000010001100110011010,
    22'b0000001101110000101001,
    22'b0000001101110000101001,
    22'b0000001111010111000011,
    22'b0000001111110101110001,
    22'b0000010001011100001010,
    22'b0000010011100001010010,
    22'b0000010001000111101100,
    22'b0000001111001100110011,
    22'b0000001101111010111000,
    22'b0000001100101000111101,
    22'b0000001011101011100001,
    22'b0000001100011110101110,
    22'b0000001101000111101100,
    22'b0000001101100110011010,
    22'b0000001110011001100110,
    22'b0000001111001100110011,
    22'b0000001111110101110001,
    22'b0000010000111101011100,
    22'b0000010010001111010111,
    22'b0000010011100001010010,
    22'b0000010100110011001101,
    22'b0000010110000101001000,
    22'b0000010111010111000011,
    22'b0000011000001010001111,
    22'b0000011000110011001101,
    22'b0000011001011100001010,
    22'b0000011001010001111011,
    22'b0000011001010001111011,
    22'b0000011000110011001101,
    22'b0000010111000010100100,
    22'b0000001111101011100001,
    22'b0000001101110000101001,
    22'b0000001011010111000011,
    22'b0000001001100110011010,
    22'b0000000111101011100001,
    22'b0000000101110000101001,
    22'b0000000011110101110001,
    22'b0000000010101110000101,
    22'b0000000010001111010111,
    22'b0000000010000101001000,
    22'b0000000010100011110110,
    22'b0000000011000010100100,
    22'b0000000011010111000011,
    22'b0000000011010111000011,
    22'b0000000011010111000011,
    22'b0000000011001100110011,
    22'b0000000010101110000101,
    22'b0000000001111010111000,
    22'b0000000001010001111011,
    22'b0000000000110011001101,
    22'b0000000000001010001111,
    22'b1111111110111000010100,
    22'b1111111110001111010111,
    22'b1111111101110000101001,
    22'b1111111101010001111011,
    22'b1111111110100011110110,
    22'b1111111110100011110110,
    22'b1111111110011001100110,
    22'b1111111110011001100110,
    22'b1111111110011001100110,
    22'b1111111110001111010111,
    22'b1111111101011100001010,
    22'b1111111100110011001101,
    22'b1111111011110101110001,
    22'b1111111010111000010100,
    22'b1111111001111010111000,
    22'b1111111001000111101100,
    22'b1111111000010100011111,
    22'b1111110111100001010010,
    22'b1111110110001111010111,
    22'b1111110100111101011100,
    22'b1111110011110101110001,
    22'b1111110001111010111000,
    22'b1111100011000010100100,
    22'b1111010111100001010010,
    22'b1111001111001100110011,
    22'b1111000111000010100100,
    22'b1110111101111010111000,
    22'b1110110110011001100110,
    22'b1110110000010100011111,
    22'b1110101100011110101110,
    22'b1110101001010001111011,
    22'b1110101000001010001111,
    22'b1110101000011110101110,
    22'b1110101001000111101100,
    22'b1110101010000101001000,
    22'b1110101010101110000101,
    22'b1110101001010001111011,
    22'b1110100111110101110001,
    22'b1110100111010111000011,
    22'b1110101001110000101001,
    22'b1110101100111101011100,
    22'b1110110100001010001111,
    22'b1110110111001100110011,
    22'b1110111001010001111011,
    22'b1110111010011001100110,
    22'b1110111010001111010111,
    22'b1110111001110000101001,
    22'b1110111001110000101001,
    22'b1110111010001111010111,
    22'b1110111100110011001101,
    22'b1110111111101011100001,
    22'b1111000011001100110011,
    22'b1111000111010111000011,
    22'b1111001110000101001000,
    22'b1111010100000000000000,
    22'b1111011010000101001000,
    22'b1111011111000010100100,
    22'b1111100010111000010100,
    22'b1111100101011100001010,
    22'b1111100111100001010010,
    22'b1111101010100011110110,
    22'b1111101101010001111011,
    22'b1111110000000000000000,
    22'b1111110010000101001000,
    22'b1111110100011110101110,
    22'b1111110110001111010111,
    22'b1111110111100001010010,
    22'b1111111011110101110001,
    22'b1111111011110101110001,
    22'b1111111011100001010010,
    22'b1111111011100001010010,
    22'b1111111011110101110001,
    22'b1111111100010100011111,
    22'b1111111100111101011100,
    22'b1111111101011100001010,
    22'b1111111110011001100110,
    22'b1111111110111000010100,
    22'b1111111111010111000011,
    22'b0000000000010100011111,
    22'b0000000001011100001010,
    22'b0000000010101110000101,
    22'b0000000100001010001111,
    22'b0000000101111010111000,
    22'b0000000111001100110011,
    22'b0000001000010100011111,
    22'b0000001001111010111000,
    22'b0000001011001100110011,
    22'b0000001100011110101110,
    22'b0000001101111010111000,
    22'b0000001111100001010010,
    22'b0000010001000111101100,
    22'b0000010000101000111101,
    22'b0000001111100001010010,
    22'b0000001110100011110110,
    22'b0000001101011100001010,
    22'b0000001100001010001111,
    22'b0000001010011001100110,
    22'b0000001001000111101100,
    22'b0000000111101011100001,
    22'b0000000100110011001101,
    22'b0000000010000101001000,
    22'b0000000000000000000000,
    22'b1111111110001111010111,
    22'b1111111100101000111101,
    22'b1111111011000010100100,
    22'b1111111010011001100110,
    22'b1111111001111010111000,
    22'b1111111011001100110011,
    22'b1111111100011110101110,
    22'b1111111101111010111000,
    22'b1111111111101011100001,
    22'b0000000011001100110011,
    22'b0000000110100011110110,
    22'b0000001001110000101001,
    22'b0000001100111101011100,
    22'b0000010000101000111101,
    22'b0000010010111000010100,
    22'b0000010010001111010111,
    22'b0000001111100001010010,
    22'b0000001110011001100110,
    22'b0000001111001100110011,
    22'b0000010001000111101100,
    22'b0000010010111000010100,
    22'b0000010010011001100110,
    22'b0000010011001100110011,
    22'b0000011111110101110001,
    22'b0000100010111000010100,
    22'b0000100101000111101100,
    22'b0000100111101011100001,
    22'b0000101000111101011100,
    22'b0000100111010111000011,
    22'b0000100101000111101100,
    22'b0000100001011100001010,
    22'b0000011101111010111000,
    22'b0000011010100011110110,
    22'b0000010100110011001101,
    22'b0000001111010111000011,
    22'b0000001010000101001000,
    22'b0000000100001010001111,
    22'b1111111111101011100001,
    22'b1111111101000111101100,
    22'b1111111001011100001010,
    22'b1111110110101110000101,
    22'b1111110100110011001101,
    22'b1111110011110101110001,
    22'b1111110010011001100110,
    22'b1111110001110000101001,
    22'b1111110001111010111000,
    22'b1111110010011001100110,
    22'b1111110010100011110110,
    22'b1111110010111000010100,
    22'b1111110011000010100100,
    22'b1111110011100001010010,
    22'b1111110011110101110001,
    22'b1111110011101011100001,
    22'b1111110011001100110011,
    22'b1111110100000000000000,
    22'b1111110100011110101110,
    22'b1111110100010100011111,
    22'b1111110100010100011111,
    22'b1111110100000000000000,
    22'b1111110011100001010010,
    22'b1111110011001100110011,
    22'b1111110010101110000101,
    22'b1111110001111010111000,
    22'b1111110000111101011100,
    22'b1111101111110101110001,
    22'b1111101110001111010111,
    22'b1111101100111101011100,
    22'b1111101011100001010010,
    22'b1111101010001111010111,
    22'b1111101000111101011100,
    22'b1111101000010100011111,
    22'b1111100111101011100001,
    22'b1111100111000010100100,
    22'b1111100110101110000101,
    22'b1111100110000101001000,
    22'b1111100101000111101100,
    22'b1111100011110101110001,
    22'b1111100010111000010100,
    22'b1111100001100110011010,
    22'b1111100000101000111101,
    22'b1111011111101011100001,
    22'b1111011111001100110011,
    22'b1111011110101110000101,
    22'b1111011110000101001000,
    22'b1111011110001111010111,
    22'b1111011110100011110110,
    22'b1111011111010111000011,
    22'b1111100101011100001010,
    22'b1111100110000101001000,
    22'b1111100110001111010111,
    22'b1111100101111010111000,
    22'b1111100101010001111011,
    22'b1111100010101110000101,
    22'b1111011110101110000101,
    22'b1111011010101110000101,
    22'b1111010101000111101100,
    22'b1111010001111010111000,
    22'b1111010000001010001111,
    22'b1111001111100001010010,
    22'b1111001111101011100001,
    22'b1111010000011110101110,
    22'b1111010001011100001010,
    22'b1111010010011001100110,
    22'b1111010011000010100100,
    22'b1111010011000010100100,
    22'b1111010010101110000101,
    22'b1111010010001111010111,
    22'b1111010001010001111011,
    22'b1111010000011110101110,
    22'b1111001111100001010010,
    22'b1111001110011001100110,
    22'b1111001101011100001010,
    22'b1111001011110101110001,
    22'b1111001001010001111011,
    22'b1111000100101000111101,
    22'b1111000000101000111101,
    22'b1110111100111101011100,
    22'b1110111010000101001000,
    22'b1110111000000000000000,
    22'b1110110111110101110001,
    22'b1110111000011110101110,
    22'b1110111001100110011010,
    22'b1110111011100001010010,
    22'b1110111100011110101110,
    22'b1110111100111101011100,
    22'b1110111100111101011100,
    22'b1110111100000000000000,
    22'b1110111010111000010100,
    22'b1110111001010001111011,
    22'b1110110001110000101001,
    22'b1110110000101000111101,
    22'b1110101111101011100001,
    22'b1110101110011001100110,
    22'b1110101101010001111011,
    22'b1110101100101000111101,
    22'b1110101100011110101110,
    22'b1110101100011110101110,
    22'b1110101101000111101100,
    22'b1110101101111010111000,
    22'b1110101111001100110011,
    22'b1110110000110011001101,
    22'b1110110011000010100100,
    22'b1110110100111101011100,
    22'b1110110111001100110011,
    22'b1110111001011100001010,
    22'b1110111100010100011111,
    22'b1110111110101110000101,
    22'b1111000000111101011100,
    22'b1111000011001100110011,
    22'b1111000110001111010111,
    22'b1111001000001010001111,
    22'b1111001001110000101001,
    22'b1111001010111000010100,
    22'b1111001100000000000000,
    22'b1111001100010100011111,
    22'b1111001100001010001111,
    22'b1111001100000000000000,
    22'b1111001011100001010010,
    22'b1111001011001100110011,
    22'b1111001010100011110110,
    22'b1111001010000101001000,
    22'b1111001001010001111011,
    22'b1111001000011110101110,
    22'b1111000111101011100001,
    22'b1111000110111000010100,
    22'b1111000110001111010111,
    22'b1111000101100110011010,
    22'b1111000101010001111011,
    22'b1111000101000111101100,
    22'b1111000101000111101100,
    22'b1111000101011100001010,
    22'b1111000101111010111000,
    22'b1111000110101110000101,
    22'b1111000111100001010010,
    22'b1111001000011110101110,
    22'b1111001001010001111011,
    22'b1111001001011100001010,
    22'b1111001001010001111011,
    22'b1111001000011110101110,
    22'b1111000111001100110011,
    22'b1111000110000101001000,
    22'b1111000100111101011100,
    22'b1111000100001010001111,
    22'b1111000011001100110011,
    22'b1111000010011001100110,
    22'b1111000001011100001010,
    22'b1111000000111101011100,
    22'b1111000000111101011100,
    22'b1111000001010001111011,
    22'b1111000001100110011010,
    22'b1111000010001111010111,
    22'b1111000010101110000101,
    22'b1111000011001100110011,
    22'b1111000011100001010010,
    22'b1111000100000000000000
};

parameter logic signed [`GYRO_WIDTH-1:0] WZ_TEST_VECTOR[`NUM_ELEMENTS] = {
    22'b1111110101010001111011,
    22'b1111110100011110101110,
    22'b1111110100001010001111,
    22'b1111110100000000000000,
    22'b1111110011101011100001,
    22'b1111110011001100110011,
    22'b1111110010100011110110,
    22'b1111110001110000101001,
    22'b1111110000110011001101,
    22'b1111101111010111000011,
    22'b1111101110001111010111,
    22'b1111101100111101011100,
    22'b1111101011101011100001,
    22'b1111101010000101001000,
    22'b1111101001000111101100,
    22'b1111101000010100011111,
    22'b1111100111101011100001,
    22'b1111100111001100110011,
    22'b1111100111010111000011,
    22'b1111100111101011100001,
    22'b1111101000010100011111,
    22'b1111101001011100001010,
    22'b1111101010001111010111,
    22'b1111101011000010100100,
    22'b1111101011110101110001,
    22'b1111101100110011001101,
    22'b1111101101011100001010,
    22'b1111101101111010111000,
    22'b1111101110011001100110,
    22'b1111101111000010100100,
    22'b1111101111010111000011,
    22'b1111101111110101110001,
    22'b1111110000001010001111,
    22'b1111110000010100011111,
    22'b1111110000010100011111,
    22'b1111110000010100011111,
    22'b1111110000010100011111,
    22'b1111110000101000111101,
    22'b1111110001000111101100,
    22'b1111110001110000101001,
    22'b1111110010101110000101,
    22'b1111110011100001010010,
    22'b1111110100001010001111,
    22'b1111110100111101011100,
    22'b1111110101111010111000,
    22'b1111110110101110000101,
    22'b1111110111100001010010,
    22'b1111111000011110101110,
    22'b1111111001110000101001,
    22'b1111111010101110000101,
    22'b1111111011101011100001,
    22'b1111111100011110101110,
    22'b1111111101110000101001,
    22'b1111111110101110000101,
    22'b1111111111100001010010,
    22'b0000000000011110101110,
    22'b0000000001000111101100,
    22'b0000000001010001111011,
    22'b0000000001011100001010,
    22'b0000000001000111101100,
    22'b0000000000110011001101,
    22'b0000000000010100011111,
    22'b1111111111101011100001,
    22'b1111111110111000010100,
    22'b1111111110111000010100,
    22'b1111111111010111000011,
    22'b0000000000000000000000,
    22'b0000000001000111101100,
    22'b0000000001111010111000,
    22'b0000000010001111010111,
    22'b0000000010001111010111,
    22'b0000000001110000101001,
    22'b0000000001010001111011,
    22'b0000000000110011001101,
    22'b0000000000011110101110,
    22'b0000000001000111101100,
    22'b0000000011000010100100,
    22'b0000000101011100001010,
    22'b0000001000010100011111,
    22'b0000001100000000000000,
    22'b0000010001010001111011,
    22'b0000010100110011001101,
    22'b0000010110011001100110,
    22'b0000010110000101001000,
    22'b0000010011000010100100,
    22'b0000001110100011110110,
    22'b0000001011000010100100,
    22'b0000001000001010001111,
    22'b0000000101000111101100,
    22'b0000000000110011001101,
    22'b1111111101110000101001,
    22'b1111111011100001010010,
    22'b1111111010100011110110,
    22'b1111111011000010100100,
    22'b1111111100010100011111,
    22'b1111111101100110011010,
    22'b1111111110101110000101,
    22'b0000000000001010001111,
    22'b0000000001011100001010,
    22'b0000000010111000010100,
    22'b0000000011110101110001,
    22'b0000000100011110101110,
    22'b0000000100111101011100,
    22'b0000000100011110101110,
    22'b0000000011110101110001,
    22'b0000000010111000010100,
    22'b0000000000110011001101,
    22'b1111111111100001010010,
    22'b1111111110100011110110,
    22'b1111111101111010111000,
    22'b1111111101110000101001,
    22'b1111111110000101001000,
    22'b1111111110001111010111,
    22'b1111111110011001100110,
    22'b1111111110100011110110,
    22'b1111111110100011110110,
    22'b1111111110101110000101,
    22'b1111111110101110000101,
    22'b1111111110111000010100,
    22'b1111111110101110000101,
    22'b1111111110101110000101,
    22'b1111111110100011110110,
    22'b1111111110111000010100,
    22'b1111111111001100110011,
    22'b1111111110111000010100,
    22'b1111111110111000010100,
    22'b1111111111001100110011,
    22'b1111111111010111000011,
    22'b0000000000000000000000,
    22'b0000000000101000111101,
    22'b0000000001010001111011,
    22'b0000000010000101001000,
    22'b0000000010101110000101,
    22'b0000000011001100110011,
    22'b0000000011100001010010,
    22'b0000000100000000000000,
    22'b0000000100001010001111,
    22'b0000000100011110101110,
    22'b0000000100101000111101,
    22'b0000000100101000111101,
    22'b0000000100101000111101,
    22'b0000000100011110101110,
    22'b0000000100000000000000,
    22'b0000000011001100110011,
    22'b0000000010001111010111,
    22'b0000000001100110011010,
    22'b0000000000110011001101,
    22'b1111111110100011110110,
    22'b1111111100010100011111,
    22'b1111111011001100110011,
    22'b1111111010011001100110,
    22'b1111111001110000101001,
    22'b1111111001100110011010,
    22'b1111111000000000000000,
    22'b1111110111101011100001,
    22'b1111110110001111010111,
    22'b1111110101000111101100,
    22'b1111110100101000111101,
    22'b1111110101010001111011,
    22'b1111110110100011110110,
    22'b1111111000101000111101,
    22'b1111111001111010111000,
    22'b1111111010011001100110,
    22'b1111111010001111010111,
    22'b1111111010000101001000,
    22'b1111111010011001100110,
    22'b1111111011100001010010,
    22'b1111111100111101011100,
    22'b1111111111010111000011,
    22'b0000000000101000111101,
    22'b0000000001011100001010,
    22'b0000000010000101001000,
    22'b0000000010011001100110,
    22'b0000000010011001100110,
    22'b0000000010011001100110,
    22'b0000000010000101001000,
    22'b0000000010100011110110,
    22'b0000000001100110011010,
    22'b0000000000011110101110,
    22'b1111111110001111010111,
    22'b1111111001100110011010,
    22'b1111110101011100001010,
    22'b1111110010001111010111,
    22'b1111110000110011001101,
    22'b1111110100001010001111,
    22'b1111110110001111010111,
    22'b1111111000101000111101,
    22'b1111111010100011110110,
    22'b1111111101100110011010,
    22'b0000000000010100011111,
    22'b0000000011110101110001,
    22'b0000001000000000000000,
    22'b0000001110011001100110,
    22'b0000010010111000010100,
    22'b0000010110011001100110,
    22'b0000011000111101011100,
    22'b0000011011001100110011,
    22'b0000011011110101110001,
    22'b0000011011110101110001,
    22'b0000011010111000010100,
    22'b0000011000110011001101,
    22'b0000011000010100011111,
    22'b0000010111001100110011,
    22'b0000010110000101001000,
    22'b0000010100010100011111,
    22'b0000010010101110000101,
    22'b0000010000111101011100,
    22'b0000010000000000000000,
    22'b0000001111001100110011,
    22'b0000001110101110000101,
    22'b0000001101111010111000,
    22'b0000001100110011001101,
    22'b0000001011101011100001,
    22'b0000001011001100110011,
    22'b0000001011101011100001,
    22'b0000001100101000111101,
    22'b0000001101110000101001,
    22'b0000001110111000010100,
    22'b0000001111001100110011,
    22'b0000001110111000010100,
    22'b0000001110000101001000,
    22'b0000001100110011001101,
    22'b0000001011101011100001,
    22'b0000001010101110000101,
    22'b0000001001110000101001,
    22'b0000001000110011001101,
    22'b0000000111001100110011,
    22'b0000000101110000101001,
    22'b0000000100000000000000,
    22'b0000000010001111010111,
    22'b1111111111110101110001,
    22'b1111111110100011110110,
    22'b1111111101100110011010,
    22'b1111111101000111101100,
    22'b1111111101010001111011,
    22'b1111111101110000101001,
    22'b1111111110101110000101,
    22'b0000000000011110101110,
    22'b0000000010001111010111,
    22'b0000000100001010001111,
    22'b0000000110000101001000,
    22'b0000001000111101011100,
    22'b0000001011001100110011,
    22'b0000001101011100001010,
    22'b0000010000000000000000,
    22'b0000010011101011100001,
    22'b0000010100110011001101,
    22'b0000010101000111101100,
    22'b0000010100000000000000,
    22'b0000010010111000010100,
    22'b0000010011101011100001,
    22'b0000010011000010100100,
    22'b0000010100010100011111,
    22'b0000010100011110101110,
    22'b0000010100110011001101,
    22'b0000010101100110011010,
    22'b0000010111100001010010,
    22'b0000011010111000010100,
    22'b0000011110111000010100,
    22'b0000100000110011001101,
    22'b0000100001111010111000,
    22'b0000100001111010111000,
    22'b0000100001000111101100,
    22'b0000100000010100011111,
    22'b0000011111110101110001,
    22'b0000011111100001010010,
    22'b0000011111101011100001,
    22'b0000011111001100110011,
    22'b0000011110011001100110,
    22'b0000011100111101011100,
    22'b0000011011100001010010,
    22'b0000011000011110101110,
    22'b0000010101111010111000,
    22'b0000010011000010100100,
    22'b0000010000010100011111,
    22'b0000001101011100001010,
    22'b0000001011100001010010,
    22'b0000001010000101001000,
    22'b0000001000010100011111,
    22'b0000000110011001100110,
    22'b0000000100110011001101,
    22'b0000000011100001010010,
    22'b0000000010011001100110,
    22'b0000000001011100001010,
    22'b0000000001010001111011,
    22'b0000000001100110011010,
    22'b0000000010000101001000,
    22'b0000000010011001100110,
    22'b0000000010000101001000,
    22'b0000000001100110011010,
    22'b0000000001010001111011,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000001000111101100,
    22'b0000000000111101011100,
    22'b0000000000011110101110,
    22'b1111111111101011100001,
    22'b1111111111001100110011,
    22'b1111111110101110000101,
    22'b1111111110100011110110,
    22'b1111111110001111010111,
    22'b1111111110001111010111,
    22'b1111111110001111010111,
    22'b1111111110000101001000,
    22'b1111111110001111010111,
    22'b1111111110100011110110,
    22'b1111111110111000010100,
    22'b1111111111010111000011,
    22'b1111111111110101110001,
    22'b0000000000000000000000,
    22'b0000000000001010001111,
    22'b0000000000010100011111,
    22'b0000000000011110101110,
    22'b0000000000101000111101,
    22'b0000000000101000111101,
    22'b0000000000011110101110,
    22'b0000000000010100011111,
    22'b0000000000000000000000,
    22'b1111111111110101110001,
    22'b1111111111101011100001,
    22'b1111111111100001010010,
    22'b1111111111010111000011,
    22'b1111111111001100110011,
    22'b1111111111000010100100,
    22'b1111111110111000010100,
    22'b1111111110111000010100,
    22'b1111111110111000010100,
    22'b1111111111000010100100,
    22'b1111111111001100110011,
    22'b1111111111010111000011,
    22'b1111111111100001010010,
    22'b1111111111101011100001,
    22'b1111111111110101110001,
    22'b0000000000000000000000,
    22'b0000000000000000000000,
    22'b0000000000000000000000,
    22'b0000000000001010001111,
    22'b0000000000000000000000,
    22'b0000000000000000000000,
    22'b0000000000000000000000,
    22'b1111111111110101110001,
    22'b1111111111101011100001,
    22'b1111111111101011100001,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111010111000011,
    22'b1111111111010111000011,
    22'b1111111111001100110011,
    22'b1111111111010111000011,
    22'b1111111111010111000011,
    22'b1111111111010111000011,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111101011100001,
    22'b1111111111101011100001,
    22'b1111111111101011100001,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111110101110001,
    22'b1111111111101011100001,
    22'b1111111111101011100001,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111010111000011,
    22'b1111111110101110000101,
    22'b1111111101111010111000,
    22'b1111111101011100001010,
    22'b1111111101111010111000,
    22'b1111111111001100110011,
    22'b0000000001011100001010,
    22'b0000000011101011100001,
    22'b0000000101000111101100,
    22'b0000000100101000111101,
    22'b0000000010101110000101,
    22'b0000000000010100011111,
    22'b1111111110011001100110,
    22'b1111111101010001111011,
    22'b1111111101100110011010,
    22'b1111111110001111010111,
    22'b1111111110111000010100,
    22'b1111111111000010100100,
    22'b1111111110101110000101,
    22'b1111111110011001100110,
    22'b1111111110001111010111,
    22'b1111111110100011110110,
    22'b1111111111000010100100,
    22'b1111111111110101110001,
    22'b0000000000010100011111,
    22'b0000000000101000111101,
    22'b0000000000101000111101,
    22'b0000000000011110101110,
    22'b0000000000010100011111,
    22'b0000000000001010001111,
    22'b0000000000001010001111,
    22'b0000000000010100011111,
    22'b0000000000011110101110,
    22'b0000000000001010001111,
    22'b0000000000000000000000,
    22'b1111111111101011100001,
    22'b1111111111010111000011,
    22'b1111111111000010100100,
    22'b1111101111101011100001,
    22'b1111100001011100001010,
    22'b1111010110001111010111,
    22'b1111011100011110101110,
    22'b1111100010000101001000,
    22'b1111011110101110000101,
    22'b1111010111100001010010,
    22'b1111010111001100110011,
    22'b1111011001011100001010,
    22'b1111011101111010111000,
    22'b1111100010000101001000,
    22'b1111100011001100110011,
    22'b1111100010101110000101,
    22'b1111100001100110011010,
    22'b1111100001010001111011,
    22'b1111100010011001100110,
    22'b1111100101110000101001,
    22'b1111101110101110000101,
    22'b1111111000000000000000,
    22'b0000000101010001111011,
    22'b0000010100111101011100,
    22'b0000100101100110011010,
    22'b0000110000111101011100,
    22'b0000110100001010001111,
    22'b0000110101000111101100,
    22'b0000110100000000000000,
    22'b0000110101000111101100,
    22'b0000110111010111000011,
    22'b0000110111100001010010,
    22'b0000110111100001010010,
    22'b0000110101100110011010,
    22'b0000101110001111010111,
    22'b0000100101111010111000,
    22'b0000011110001111010111,
    22'b0000010110100011110110,
    22'b0000001101000111101100,
    22'b0000001000001010001111,
    22'b0000000100010100011111,
    22'b0000000000001010001111,
    22'b1111111011100001010010,
    22'b1111111000001010001111,
    22'b1111110101110000101001,
    22'b1111110101010001111011,
    22'b1111110111001100110011,
    22'b1111111010000101001000,
    22'b1111111101100110011010,
    22'b0000000010000101001000,
    22'b0000000101000111101100,
    22'b0000001000000000000000,
    22'b0000001011000010100100,
    22'b0000001110001111010111,
    22'b0000010001000111101100,
    22'b0000010010101110000101,
    22'b0000001111001100110011,
    22'b0000001011010111000011,
    22'b0000000100011110101110,
    22'b0000000001000111101100,
    22'b1111111111001100110011,
    22'b1111111110101110000101,
    22'b1111111101011100001010,
    22'b1111111100010100011111,
    22'b1111111010001111010111,
    22'b1111110111110101110001,
    22'b1111110101010001111011,
    22'b1111110100111101011100,
    22'b1111110101010001111011,
    22'b1111110110001111010111,
    22'b1111111000001010001111,
    22'b1111111001011100001010,
    22'b1111111010111000010100,
    22'b1111111100101000111101,
    22'b1111111110101110000101,
    22'b0000000000101000111101,
    22'b0000000010011001100110,
    22'b0000000100001010001111,
    22'b0000000101111010111000,
    22'b0000000110100011110110,
    22'b0000000101011100001010,
    22'b0000000100001010001111,
    22'b0000000010001111010111,
    22'b0000000001000111101100,
    22'b0000000000110011001101,
    22'b0000000000101000111101,
    22'b0000000000010100011111,
    22'b1111111111010111000011,
    22'b1111111110011001100110,
    22'b1111111101010001111011,
    22'b1111111100011110101110,
    22'b1111111100001010001111,
    22'b1111111100001010001111,
    22'b1111111100101000111101,
    22'b1111111101000111101100,
    22'b1111111101111010111000,
    22'b1111111110100011110110,
    22'b1111111111000010100100,
    22'b1111111111110101110001,
    22'b0000000000011110101110,
    22'b0000000001000111101100,
    22'b0000000001111010111000,
    22'b0000000010101110000101,
    22'b0000000010101110000101,
    22'b0000000010001111010111,
    22'b0000000001011100001010,
    22'b0000000000110011001101,
    22'b0000000000011110101110,
    22'b0000000000101000111101,
    22'b0000000000111101011100,
    22'b0000000000101000111101,
    22'b1111111111010111000011,
    22'b1111111101010001111011,
    22'b1111111100011110101110,
    22'b1111111110000101001000,
    22'b1111110101010001111011,
    22'b1111100111100001010010,
    22'b1111011110011001100110,
    22'b1111010101011100001010,
    22'b1111100100101000111101,
    22'b1111101101110000101001,
    22'b1111110010000101001000,
    22'b1111101111101011100001,
    22'b1111101110101110000101,
    22'b1111110010111000010100,
    22'b1111110111110101110001,
    22'b1111111100011110101110,
    22'b1111111111001100110011,
    22'b1111111111000010100100,
    22'b1111111100010100011111,
    22'b1111111000110011001101,
    22'b1111110100110011001101,
    22'b1111110011100001010010,
    22'b1111110100110011001101,
    22'b1111110101011100001010,
    22'b1111110100001010001111,
    22'b1111110101100110011010,
    22'b1111111101000111101100,
    22'b0000001001111010111000,
    22'b0000011011101011100001,
    22'b0000100100000000000000,
    22'b0000100101100110011010,
    22'b0000100000011110101110,
    22'b0000010100111101011100,
    22'b0000001110000101001000,
    22'b0000001011010111000011,
    22'b0000001101010001111011,
    22'b0000010001100110011010,
    22'b0000010110101110000101,
    22'b0000010111110101110001,
    22'b0000010110001111010111,
    22'b0000010011000010100100,
    22'b0000001110101110000101,
    22'b0000001100101000111101,
    22'b0000001011100001010010,
    22'b0000001100000000000000,
    22'b0000001101110000101001,
    22'b0000010000101000111101,
    22'b0000010010100011110110,
    22'b0000010011101011100001,
    22'b0000010100010100011111,
    22'b0000010100110011001101,
    22'b0000010101110000101001,
    22'b0000010111100001010010,
    22'b0000011001110000101001,
    22'b0000011011100001010010,
    22'b0000011110011001100110,
    22'b0000100000111101011100,
    22'b0000100011100001010010,
    22'b0000100101100110011010,
    22'b0000100110011001100110,
    22'b0000100110001111010111,
    22'b0000100101110000101001,
    22'b0000100100110011001101,
    22'b0000100011101011100001,
    22'b0000100010000101001000,
    22'b0000100001000111101100,
    22'b0000100000000000000000,
    22'b0000011111100001010010,
    22'b0000011111100001010010,
    22'b0000100000000000000000,
    22'b0000100000010100011111,
    22'b0000100000000000000000,
    22'b0000011111001100110011,
    22'b0000011101011100001010,
    22'b0000011100011110101110,
    22'b0000011100000000000000,
    22'b0000011011101011100001,
    22'b0000011011101011100001,
    22'b0000011011000010100100,
    22'b0000010100111101011100,
    22'b0000001100011110101110,
    22'b0000000010100011110110,
    22'b1111111111110101110001,
    22'b0000000001111010111000,
    22'b0000001000000000000000,
    22'b0000001111010111000011,
    22'b0000010111001100110011,
    22'b0000011100001010001111,
    22'b0000100000101000111101,
    22'b0000100100101000111101,
    22'b0000101001000111101100,
    22'b0000101100011110101110,
    22'b0000101110001111010111,
    22'b0000101101111010111000,
    22'b0000101101111010111000,
    22'b0000101100010100011111,
    22'b0000101101111010111000,
    22'b0000110001111010111000,
    22'b0000110110111000010100,
    22'b0000111011100001010010,
    22'b0000111100010100011111,
    22'b0000111010011001100110,
    22'b0000110111100001010010,
    22'b0000110010011001100110,
    22'b0000101110101110000101,
    22'b0000101010101110000101,
    22'b0000100111010111000011,
    22'b0000100010011001100110,
    22'b0000011110001111010111,
    22'b0000011001111010111000,
    22'b0000010101110000101001,
    22'b0000001100000000000000,
    22'b0000000001100110011010,
    22'b1111110011100001010010,
    22'b1111100010001111010111,
    22'b1111001010011001100110,
    22'b1110110111001100110011,
    22'b1110110001110000101001,
    22'b1111001000000000000000,
    22'b1111011100101000111101,
    22'b1111110010100011110110,
    22'b0000001000111101011100,
    22'b0000011100110011001101,
    22'b0000101100101000111101,
    22'b0000101111100001010010,
    22'b0000101100110011001101,
    22'b0000100101100110011010,
    22'b0000011100010100011111,
    22'b0000010000011110101110,
    22'b0000001001111010111000,
    22'b0000000111001100110011,
    22'b0000000110011001100110,
    22'b0000000101000111101100,
    22'b0000000011101011100001,
    22'b0000000010000101001000,
    22'b0000000000101000111101,
    22'b1111111111000010100100,
    22'b1111111110001111010111,
    22'b1111111111100001010010,
    22'b0000000010000101001000,
    22'b0000000101110000101001,
    22'b0000001010001111010111,
    22'b0000001101110000101001,
    22'b0000010000010100011111,
    22'b0000010010100011110110,
    22'b0000010100001010001111,
    22'b0000010011010111000011,
    22'b0000010001110000101001,
    22'b0000001111100001010010,
    22'b0000001101000111101100,
    22'b0000001001111010111000,
    22'b0000001001000111101100,
    22'b0000001001011100001010,
    22'b0000001010111000010100,
    22'b0000001100010100011111,
    22'b0000001101011100001010,
    22'b0000001100111101011100,
    22'b0000001100011110101110,
    22'b0000001100001010001111,
    22'b0000001100010100011111,
    22'b0000001100001010001111,
    22'b0000001011001100110011,
    22'b0000001000111101011100,
    22'b0000000100000000000000,
    22'b1111111111000010100100,
    22'b1111111001011100001010,
    22'b1111110011010111000011,
    22'b1111101101010001111011,
    22'b1111100101000111101100,
    22'b1111011111100001010010,
    22'b1111011010111000010100,
    22'b1111010110101110000101,
    22'b1111010010001111010111,
    22'b1111010000000000000000,
    22'b1111001110111000010100,
    22'b1111001111000010100100,
    22'b1111010001010001111011,
    22'b1111010100110011001101,
    22'b1111011001011100001010,
    22'b1111011111001100110011,
    22'b1111100111110101110001,
    22'b1111101111001100110011,
    22'b1111110110000101001000,
    22'b1111111011101011100001,
    22'b0000000000111101011100,
    22'b0000000011010111000011,
    22'b0000000100101000111101,
    22'b0000000100111101011100,
    22'b0000000100110011001101,
    22'b0000000100011110101110,
    22'b0000000100010100011111,
    22'b0000000100000000000000,
    22'b0000000011100001010010,
    22'b0000000010100011110110,
    22'b0000000001100110011010,
    22'b0000000000110011001101,
    22'b1111111111110101110001,
    22'b1111111111000010100100,
    22'b1111111101110000101001,
    22'b1111111100110011001101,
    22'b1111111100000000000000,
    22'b1111111011010111000011,
    22'b1111111010011001100110,
    22'b1111111001011100001010,
    22'b1111111000011110101110,
    22'b1111110111000010100100,
    22'b1111110100001010001111,
    22'b1111110001000111101100,
    22'b1111101110000101001000,
    22'b1111101001010001111011,
    22'b1111100101110000101001,
    22'b1111100010011001100110,
    22'b1111011111010111000011,
    22'b1111011011110101110001,
    22'b1111011010100011110110,
    22'b1111011001100110011010,
    22'b1111011000111101011100,
    22'b1111011000010100011111,
    22'b1111010111101011100001,
    22'b1111011010111000010100,
    22'b1111011100111101011100,
    22'b1111100010001111010111,
    22'b1111100110111000010100,
    22'b1111101011101011100001,
    22'b1111101110111000010100,
    22'b1111110000101000111101,
    22'b1111110000101000111101,
    22'b1111101110111000010100,
    22'b1111101100000000000000,
    22'b1111101010111000010100,
    22'b1111101010101110000101,
    22'b1111101011001100110011,
    22'b1111101100001010001111,
    22'b1111101100101000111101,
    22'b1111101101010001111011,
    22'b1111101110000101001000,
    22'b1111101110101110000101,
    22'b1111101110111000010100,
    22'b1111101111000010100100,
    22'b1111101111010111000011,
    22'b1111110000000000000000,
    22'b1111110001000111101100,
    22'b1111110010100011110110,
    22'b1111110100010100011111,
    22'b1111110111000010100100,
    22'b1111111001011100001010,
    22'b1111111011101011100001,
    22'b1111111110000101001000,
    22'b0000000000010100011111,
    22'b0000000010111000010100,
    22'b0000000101000111101100,
    22'b0000001000111101011100,
    22'b0000001100001010001111,
    22'b0000001111000010100100,
    22'b0000010001100110011010,
    22'b0000010100000000000000,
    22'b0000010110111000010100,
    22'b0000011000011110101110,
    22'b0000011001111010111000,
    22'b0000011011101011100001,
    22'b0000011101000111101100,
    22'b0000011110011001100110,
    22'b0000011111110101110001,
    22'b0000100001110000101001,
    22'b0000100011100001010010,
    22'b0000100101010001111011,
    22'b0000100101010001111011,
    22'b0000100100011110101110,
    22'b0000100010111000010100,
    22'b0000100000111101011100,
    22'b0000100000110011001101,
    22'b0000100010111000010100,
    22'b0000100110111000010100,
    22'b0000101101010001111011,
    22'b0000110101100110011010,
    22'b0000110101000111101100,
    22'b0000101101111010111000,
    22'b0000100100011110101110,
    22'b0000011011000010100100,
    22'b0000001111001100110011,
    22'b0000000111100001010010,
    22'b0000000010100011110110,
    22'b0000000001010001111011,
    22'b0000000011010111000011,
    22'b0000000101110000101001,
    22'b0000000111101011100001,
    22'b0000001001011100001010,
    22'b0000001010111000010100,
    22'b0000001100101000111101,
    22'b0000001101110000101001,
    22'b0000001111001100110011,
    22'b0000010000111101011100,
    22'b0000010011100001010010,
    22'b0000010101100110011010,
    22'b0000010111010111000011,
    22'b0000011000101000111101,
    22'b0000011001100110011010,
    22'b0000011001010001111011,
    22'b0000011000010100011111,
    22'b0000010111001100110011,
    22'b0000010101100110011010,
    22'b0000010100110011001101,
    22'b0000010100101000111101,
    22'b0000010100000000000000,
    22'b0000010011100001010010,
    22'b0000010100110011001101,
    22'b0000010101000111101100,
    22'b0000010101100110011010,
    22'b0000010110011001100110,
    22'b0000010110100011110110,
    22'b0000010110001111010111,
    22'b0000010101111010111000,
    22'b0000010101100110011010,
    22'b0000010101011100001010,
    22'b0000010101111010111000,
    22'b0000010110001111010111,
    22'b0000010110111000010100,
    22'b0000010111101011100001,
    22'b0000011000110011001101,
    22'b0000011001111010111000,
    22'b0000011011000010100100,
    22'b0000011100001010001111,
    22'b0000011100111101011100,
    22'b0000011101011100001010,
    22'b0000011101110000101001,
    22'b0000011110011001100110,
    22'b0000011111001100110011,
    22'b0000100000011110101110,
    22'b0000100001010001111011,
    22'b0000100001111010111000,
    22'b0000100010000101001000,
    22'b0000100001111010111000,
    22'b0000100000111101011100,
    22'b0000011111110101110001,
    22'b0000011110001111010111,
    22'b0000011100101000111101,
    22'b0000011010100011110110,
    22'b0000011000111101011100,
    22'b0000010111101011100001,
    22'b0000010110100011110110,
    22'b0000010101010001111011,
    22'b0000010100011110101110,
    22'b0000010011100001010010,
    22'b0000010010111000010100,
    22'b0000010010000101001000,
    22'b0000010001011100001010,
    22'b0000010000111101011100,
    22'b0000010000010100011111,
    22'b0000001111110101110001,
    22'b0000001111101011100001,
    22'b0000001111101011100001,
    22'b0000001111100001010010,
    22'b0000001111101011100001,
    22'b0000001111101011100001,
    22'b0000001111101011100001,
    22'b0000001111101011100001,
    22'b0000001111100001010010,
    22'b0000001111000010100100,
    22'b0000001110011001100110,
    22'b0000001101100110011010,
    22'b0000001100101000111101,
    22'b0000001011100001010010,
    22'b0000001010000101001000,
    22'b0000001000111101011100,
    22'b0000000111110101110001,
    22'b0000000110001111010111,
    22'b0000000100000000000000,
    22'b0000000011001100110011,
    22'b0000000001011100001010,
    22'b1111111111001100110011,
    22'b1111111100011110101110,
    22'b1111111011000010100100,
    22'b1111111001111010111000,
    22'b1111111000011110101110,
    22'b1111110111100001010010,
    22'b1111110111000010100100,
    22'b1111110110100011110110,
    22'b1111110110100011110110,
    22'b1111110101100110011010,
    22'b1111110101000111101100,
    22'b1111110100111101011100,
    22'b1111110100111101011100,
    22'b1111110100011110101110,
    22'b1111110011100001010010,
    22'b1111110001111010111000,
    22'b1111110000010100011111,
    22'b1111101110011001100110,
    22'b1111101010101110000101,
    22'b1111101000001010001111,
    22'b1111100100111101011100,
    22'b1111100010100011110110,
    22'b1111100010011001100110,
    22'b1111100011100001010010,
    22'b1111100101111010111000,
    22'b1111101001010001111011,
    22'b1111110001000111101100,
    22'b1111111010100011110110,
    22'b0000000110001111010111,
    22'b0000010010101110000101,
    22'b0000011011101011100001,
    22'b0000011011000010100100,
    22'b0000011001011100001010,
    22'b0000011010111000010100,
    22'b0000100000111101011100,
    22'b0000110000001010001111,
    22'b0000111010001111010111,
    22'b0000111110101110000101,
    22'b0001000010001111010111,
    22'b0001000100010100011111,
    22'b0000111110100011110110,
    22'b0000110101010001111011,
    22'b0000101100111101011100,
    22'b0000100110101110000101,
    22'b0000100000111101011100,
    22'b0000011100000000000000,
    22'b0000011000001010001111,
    22'b0000010100010100011111,
    22'b0000001110100011110110,
    22'b0000001010111000010100,
    22'b0000000111110101110001,
    22'b0000000101010001111011,
    22'b0000000001110000101001,
    22'b1111110100010100011111,
    22'b1111110001100110011010,
    22'b1111101111110101110001,
    22'b1111110000011110101110,
    22'b1111110011101011100001,
    22'b1111111001011100001010,
    22'b1111111111001100110011,
    22'b0000000110001111010111,
    22'b0000001100001010001111,
    22'b0000010001111010111000,
    22'b0000010110111000010100,
    22'b0000011011110101110001,
    22'b0000011100000000000000,
    22'b0000011000011110101110,
    22'b0000010010111000010100,
    22'b0000001001110000101001,
    22'b0000000101011100001010,
    22'b0000000001011100001010,
    22'b1111111100011110101110,
    22'b1111111000110011001101,
    22'b1111110111110101110001,
    22'b1111110110000101001000,
    22'b1111110001111010111000,
    22'b1111110101111010111000,
    22'b1111111010011001100110,
    22'b1111111011010111000011,
    22'b1111111011000010100100,
    22'b1111111100001010001111,
    22'b1111111101111010111000,
    22'b0000000000000000000000,
    22'b0000000001010001111011,
    22'b0000000000111101011100,
    22'b0000000001100110011010,
    22'b0000000011000010100100,
    22'b0000000100001010001111,
    22'b0000000100011110101110,
    22'b0000000010101110000101,
    22'b1111111111010111000011,
    22'b1111111010100011110110,
    22'b1111110111001100110011,
    22'b1111110011110101110001,
    22'b1111110000010100011111,
    22'b1111101101100110011010,
    22'b1111101010101110000101,
    22'b1111101100010100011111,
    22'b1111101111000010100100,
    22'b1111110000001010001111,
    22'b1111101111101011100001,
    22'b1111110000011110101110,
    22'b1111110010000101001000,
    22'b1111110011001100110011,
    22'b1111110011010111000011,
    22'b1111110011001100110011,
    22'b1111110011100001010010,
    22'b1111110100000000000000,
    22'b1111110100011110101110,
    22'b1111110100101000111101,
    22'b1111110101100110011010,
    22'b1111110111110101110001,
    22'b0000000100000000000000,
    22'b0000000111101011100001,
    22'b0000001001110000101001,
    22'b0000001011001100110011,
    22'b0000001011101011100001,
    22'b0000001011010111000011,
    22'b0000001001010001111011,
    22'b0000000110101110000101,
    22'b0000000011101011100001,
    22'b0000000000011110101110,
    22'b1111111100000000000000,
    22'b1111111001000111101100,
    22'b1111110110100011110110,
    22'b1111110100001010001111,
    22'b1111110000110011001101,
    22'b1111101110100011110110,
    22'b1111101100111101011100,
    22'b1111101011110101110001,
    22'b1111101011001100110011,
    22'b1111101011010111000011,
    22'b1111101011110101110001,
    22'b1111101100010100011111,
    22'b1111101101000111101100,
    22'b1111101101111010111000,
    22'b1111101101111010111000,
    22'b1111101110011001100110,
    22'b1111101110001111010111,
    22'b1111101110011001100110,
    22'b1111101110100011110110,
    22'b1111101111010111000011,
    22'b1111110000010100011111,
    22'b1111110001111010111000,
    22'b1111110100000000000000,
    22'b1111110110000101001000,
    22'b1111111000000000000000,
    22'b1111111010000101001000,
    22'b1111111100001010001111,
    22'b1111111111001100110011,
    22'b0000000001100110011010,
    22'b0000000100001010001111,
    22'b0000000111010111000011,
    22'b0000001100000000000000,
    22'b0000001111000010100100,
    22'b0000010011010111000011,
    22'b0000010111010111000011,
    22'b0000011100101000111101,
    22'b0000100001110000101001,
    22'b0000100101100110011010,
    22'b0000101010000101001000,
    22'b0000101100110011001101,
    22'b0000110010000101001000,
    22'b0000110011110101110001,
    22'b0000110101111010111000,
    22'b0000110110101110000101,
    22'b0000111000110011001101,
    22'b0000111000101000111101,
    22'b0000111010011001100110,
    22'b0000111010111000010100,
    22'b0000111010111000010100,
    22'b0000111011101011100001,
    22'b0000111100000000000000,
    22'b0000111011110101110001,
    22'b0000111010101110000101,
    22'b0000111010011001100110,
    22'b0000111001100110011010,
    22'b0000111001000111101100,
    22'b0000111000011110101110,
    22'b0000110110001111010111,
    22'b0000110011110101110001,
    22'b0000110001010001111011,
    22'b0000101110101110000101,
    22'b0000101101100110011010,
    22'b0000101101000111101100,
    22'b0000101100000000000000,
    22'b0000101010101110000101,
    22'b0000101000111101011100,
    22'b0000100110100011110110,
    22'b0000100101011100001010,
    22'b0000100100011110101110,
    22'b0000100101011100001010,
    22'b0000100110011001100110,
    22'b0000100100011110101110,
    22'b0000100010100011110110,
    22'b0000100000010100011111,
    22'b0000011101011100001010,
    22'b0000011010000101001000,
    22'b0000010100111101011100,
    22'b0000010001110000101001,
    22'b0000001111001100110011,
    22'b0000001100000000000000,
    22'b0000000111001100110011,
    22'b0000000011101011100001,
    22'b1111111111110101110001,
    22'b1111111011100001010010,
    22'b1111110111001100110011,
    22'b1111110000101000111101,
    22'b1111101100001010001111,
    22'b1111100110111000010100,
    22'b1111100010011001100110,
    22'b1111011010100011110110,
    22'b1111010110101110000101,
    22'b1111010111000010100100,
    22'b1111011000101000111101,
    22'b1111011010001111010111,
    22'b1111100000000000000000,
    22'b1111100100010100011111,
    22'b1111100111110101110001,
    22'b1111101001100110011010,
    22'b1111101001110000101001,
    22'b1111101000111101011100,
    22'b1111100111101011100001,
    22'b1111100100111101011100,
    22'b1111011110101110000101,
    22'b1111011100001010001111,
    22'b1111011000110011001101,
    22'b1111010110011001100110,
    22'b1111010111100001010010,
    22'b1111011000110011001101,
    22'b1111011000110011001101,
    22'b1111010111110101110001,
    22'b1111010111110101110001,
    22'b1111011001111010111000,
    22'b1111011011010111000011,
    22'b1111011011101011100001,
    22'b1111011010100011110110,
    22'b1111010110101110000101,
    22'b1111001110111000010100,
    22'b1111000111010111000011,
    22'b1111000100000000000000,
    22'b1111000100101000111101,
    22'b1111000111100001010010,
    22'b1111001110011001100110,
    22'b1111010101000111101100,
    22'b1111011010100011110110,
    22'b1111011101000111101100,
    22'b1111011111001100110011,
    22'b1111100000111101011100,
    22'b1111100011101011100001,
    22'b1111100101110000101001,
    22'b1111100111101011100001,
    22'b1111101001000111101100,
    22'b1111101010011001100110,
    22'b1111101011001100110011,
    22'b1111101011110101110001,
    22'b1111101100010100011111,
    22'b1111101100010100011111,
    22'b1111101100001010001111,
    22'b1111101011110101110001,
    22'b1111101011000010100100,
    22'b1111101000101000111101,
    22'b1111100010001111010111,
    22'b1111011011001100110011,
    22'b1111010101110000101001,
    22'b1111010011000010100100,
    22'b1111010100000000000000,
    22'b1111010111010111000011,
    22'b1111011100010100011111,
    22'b1111100001011100001010,
    22'b1111100101100110011010,
    22'b1111100101011100001010,
    22'b1111100101111010111000,
    22'b1111100101110000101001,
    22'b1111100100101000111101,
    22'b1111100100010100011111,
    22'b1111100011100001010010,
    22'b1111100011101011100001,
    22'b1111100101111010111000,
    22'b1111101001000111101100,
    22'b1111101100011110101110,
    22'b1111110000001010001111,
    22'b1111110101100110011010,
    22'b1111111001011100001010,
    22'b1111111100001010001111,
    22'b1111111110001111010111,
    22'b0000000001000111101100,
    22'b0000000000101000111101,
    22'b1111111110111000010100,
    22'b1111111010111000010100,
    22'b1111110100011110101110,
    22'b1111100110011001100110,
    22'b1111010000101000111101,
    22'b1111000100110011001101,
    22'b1110111100001010001111,
    22'b1110111001000111101100,
    22'b1110111100011110101110,
    22'b1111000011001100110011,
    22'b1111001010011001100110,
    22'b1111010001010001111011,
    22'b1111011001010001111011,
    22'b1111011110101110000101,
    22'b1111100011010111000011,
    22'b1111100111101011100001,
    22'b1111101100001010001111,
    22'b1111101101111010111000,
    22'b1111101110001111010111,
    22'b1111101100110011001101,
    22'b1111101010100011110110,
    22'b1111101000001010001111,
    22'b1111100110001111010111,
    22'b1111100100111101011100,
    22'b1111100100011110101110,
    22'b1111100100011110101110,
    22'b1111100100011110101110,
    22'b1111100110011001100110,
    22'b1111101010101110000101,
    22'b1111101111110101110001,
    22'b1111110100000000000000,
    22'b1111110110011001100110,
    22'b1111110101000111101100,
    22'b1111110011010111000011,
    22'b1111110001110000101001,
    22'b1111101111101011100001,
    22'b1111101101110000101001,
    22'b1111101011100001010010,
    22'b1111100111010111000011,
    22'b1111100000001010001111,
    22'b1111011101000111101100,
    22'b1111011011010111000011,
    22'b1111011001010001111011,
    22'b1111011000010100011111,
    22'b1111011010000101001000,
    22'b1111011100011110101110,
    22'b1111011110100011110110,
    22'b1111100000011110101110,
    22'b1111100001010001111011,
    22'b1111100001111010111000,
    22'b1111100010100011110110,
    22'b1111100010011001100110,
    22'b1111100010100011110110,
    22'b1111100100010100011111,
    22'b1111100101110000101001,
    22'b1111100110000101001000,
    22'b1111100110001111010111,
    22'b1111100110111000010100,
    22'b1111101000000000000000,
    22'b1111101001111010111000,
    22'b1111101011010111000011,
    22'b1111101100011110101110,
    22'b1111101101010001111011,
    22'b1111101101010001111011,
    22'b1111101100111101011100,
    22'b1111101100011110101110,
    22'b1111101100000000000000,
    22'b1111101011101011100001,
    22'b1111101011001100110011,
    22'b1111101011000010100100,
    22'b1111101011000010100100,
    22'b1111101010111000010100,
    22'b1111101010100011110110,
    22'b1111101010000101001000,
    22'b1111101001100110011010,
    22'b1111101001000111101100,
    22'b1111101000110011001101,
    22'b1111101000001010001111,
    22'b1111100111100001010010,
    22'b1111100110100011110110,
    22'b1111100101100110011010,
    22'b1111100100000000000000,
    22'b1111100010111000010100,
    22'b1111100001111010111000,
    22'b1111100001000111101100,
    22'b1111100000101000111101,
    22'b1111100000101000111101,
    22'b1111100000101000111101,
    22'b1111100000111101011100,
    22'b1111100001010001111011,
    22'b1111100010001111010111,
    22'b1111100011100001010010,
    22'b1111100100111101011100,
    22'b1111100110101110000101,
    22'b1111101001000111101100,
    22'b1111101010101110000101,
    22'b1111101011101011100001,
    22'b1111101011001100110011,
    22'b1111101010100011110110,
    22'b1111101010100011110110,
    22'b1111101011000010100100,
    22'b1111101010111000010100,
    22'b1111101010001111010111,
    22'b1111101001110000101001,
    22'b1111101001010001111011,
    22'b1111101000101000111101,
    22'b1111101000010100011111,
    22'b1111100111110101110001,
    22'b1111100110111000010100,
    22'b1111100100101000111101,
    22'b1111100001111010111000,
    22'b1111011110100011110110,
    22'b1111011010100011110110,
    22'b1111010100011110101110,
    22'b1111001111100001010010,
    22'b1111001011001100110011,
    22'b1111001000001010001111,
    22'b1111000110011001100110,
    22'b1111000110011001100110,
    22'b1111000110111000010100,
    22'b1111000111100001010010,
    22'b1111001000110011001101,
    22'b1111001001110000101001,
    22'b1111001011000010100100,
    22'b1111001101010001111011,
    22'b1111010010001111010111,
    22'b1111010111010111000011,
    22'b1111011100111101011100,
    22'b1111100001111010111000,
    22'b1111100101110000101001,
    22'b1111101001010001111011,
    22'b1111101011010111000011,
    22'b1111101101010001111011,
    22'b1111101111010111000011,
    22'b1111110010000101001000,
    22'b1111110100001010001111,
    22'b1111110110100011110110,
    22'b1111111001111010111000,
    22'b1111111100011110101110,
    22'b1111111110111000010100,
    22'b0000000000101000111101,
    22'b0000000001111010111000,
    22'b0000000010100011110110,
    22'b0000000010111000010100,
    22'b0000000010101110000101,
    22'b0000000010100011110110,
    22'b0000000010100011110110,
    22'b0000000010011001100110,
    22'b0000000010011001100110,
    22'b0000000010011001100110,
    22'b0000000010011001100110,
    22'b0000000010001111010111,
    22'b0000000010000101001000,
    22'b0000000001111010111000,
    22'b0000000001011100001010,
    22'b0000000001000111101100,
    22'b0000000000111101011100,
    22'b0000000000110011001101,
    22'b0000000000110011001101,
    22'b0000000001000111101100,
    22'b0000000001011100001010,
    22'b0000000010000101001000,
    22'b0000000011000010100100,
    22'b0000000100001010001111,
    22'b0000000101000111101100,
    22'b0000000110000101001000,
    22'b0000000110111000010100,
    22'b0000000111101011100001,
    22'b0000001000011110101110,
    22'b0000001001010001111011,
    22'b0000001010001111010111,
    22'b0000001011001100110011,
    22'b0000001100111101011100,
    22'b0000001110100011110110,
    22'b0000010000001010001111,
    22'b0000010001000111101100,
    22'b0000010010011001100110,
    22'b0000010011010111000011,
    22'b0000010100000000000000,
    22'b0000010101110000101001,
    22'b0000011000101000111101,
    22'b0000011101111010111000,
    22'b0000011111110101110001,
    22'b0000100000111101011100,
    22'b0000100001011100001010,
    22'b0000100001110000101001,
    22'b0000100010100011110110,
    22'b0000100011001100110011,
    22'b0000100011101011100001,
    22'b0000100011110101110001,
    22'b0000100101010001111011,
    22'b0000100101011100001010,
    22'b0000100101010001111011,
    22'b0000100110000101001000,
    22'b0000100110101110000101,
    22'b0000100110111000010100,
    22'b0000100111001100110011,
    22'b0000100111110101110001,
    22'b0000101000001010001111,
    22'b0000101000011110101110,
    22'b0000101000011110101110,
    22'b0000101000000000000000,
    22'b0000100111001100110011,
    22'b0000100110001111010111,
    22'b0000100011101011100001,
    22'b0000100001100110011010,
    22'b0000011110101110000101,
    22'b0000011110000101001000,
    22'b0000100000011110101110,
    22'b0000100110011001100110,
    22'b0000100111110101110001,
    22'b0000100100101000111101,
    22'b0000100000101000111101,
    22'b0000011110001111010111,
    22'b0000011011100001010010,
    22'b0000011000101000111101,
    22'b0000010100111101011100,
    22'b0000010001110000101001,
    22'b0000001111000010100100,
    22'b0000001111110101110001,
    22'b0000010001100110011010,
    22'b0000010011000010100100,
    22'b0000010100001010001111,
    22'b0000010100001010001111,
    22'b0000010011110101110001,
    22'b0000010010111000010100,
    22'b0000010001110000101001,
    22'b0000010000001010001111,
    22'b0000001110100011110110,
    22'b0000001110011001100110,
    22'b0000001110100011110110,
    22'b0000001111000010100100,
    22'b0000001111101011100001,
    22'b0000010000001010001111,
    22'b0000010000101000111101,
    22'b0000010000111101011100,
    22'b0000010001011100001010,
    22'b0000010001000111101100,
    22'b0000001110111000010100,
    22'b0000001100110011001101,
    22'b0000001100111101011100,
    22'b0000001010100011110110,
    22'b0000001011001100110011,
    22'b0000001010100011110110,
    22'b0000001001100110011010,
    22'b0000001000101000111101,
    22'b0000001000000000000000,
    22'b0000001000010100011111,
    22'b0000001001011100001010,
    22'b0000001011110101110001,
    22'b0000001101010001111011,
    22'b0000001111100001010010,
    22'b0000010000001010001111,
    22'b0000001111010111000011,
    22'b0000001100011110101110,
    22'b0000001010000101001000,
    22'b0000000110001111010111,
    22'b0000000100000000000000,
    22'b0000000010111000010100,
    22'b0000000010101110000101,
    22'b0000000011000010100100,
    22'b0000000011010111000011,
    22'b0000000011100001010010,
    22'b0000000011001100110011,
    22'b0000000010111000010100,
    22'b0000000010101110000101,
    22'b0000000010111000010100,
    22'b0000000011001100110011,
    22'b0000000011101011100001,
    22'b0000000100010100011111,
    22'b0000000100111101011100,
    22'b0000000101100110011010,
    22'b0000000110000101001000,
    22'b0000000110001111010111,
    22'b0000000110001111010111,
    22'b0000000110011001100110,
    22'b0000000110011001100110,
    22'b0000000110101110000101,
    22'b0000000111000010100100,
    22'b0000000111100001010010,
    22'b0000001000000000000000,
    22'b0000001000110011001101,
    22'b0000001001000111101100,
    22'b0000001001000111101100,
    22'b0000001000110011001101,
    22'b0000001000010100011111,
    22'b0000001000000000000000,
    22'b0000001000000000000000,
    22'b0000001000000000000000,
    22'b0000001000001010001111,
    22'b0000001000001010001111,
    22'b0000001000010100011111,
    22'b0000001000011110101110,
    22'b0000001000110011001101,
    22'b0000001001010001111011,
    22'b0000001001100110011010,
    22'b0000001001110000101001,
    22'b0000001001110000101001,
    22'b0000001001100110011010,
    22'b0000001001000111101100,
    22'b0000001000101000111101,
    22'b0000000111010111000011,
    22'b0000001000000000000000,
    22'b0000001010001111010111,
    22'b0000001100011110101110,
    22'b0000001110111000010100,
    22'b0000010000101000111101,
    22'b0000010001100110011010,
    22'b0000010010101110000101,
    22'b0000010010101110000101,
    22'b0000010001011100001010,
    22'b0000010000001010001111,
    22'b0000001110101110000101,
    22'b0000001101010001111011,
    22'b0000001011001100110011,
    22'b0000001001100110011010,
    22'b0000001000001010001111,
    22'b0000000111001100110011,
    22'b0000000110100011110110,
    22'b0000000110000101001000,
    22'b0000000101111010111000,
    22'b0000000110000101001000,
    22'b0000000110111000010100,
    22'b0000000111110101110001,
    22'b0000001000101000111101,
    22'b0000001001010001111011,
    22'b0000001001111010111000,
    22'b0000001010011001100110,
    22'b0000001010101110000101,
    22'b0000001010111000010100,
    22'b0000001011000010100100,
    22'b0000001011000010100100,
    22'b0000001010111000010100,
    22'b0000001010000101001000,
    22'b0000001001010001111011,
    22'b0000001000010100011111,
    22'b0000000111001100110011,
    22'b0000000110000101001000,
    22'b0000000100111101011100,
    22'b0000000100011110101110,
    22'b0000000100011110101110,
    22'b0000000100110011001101,
    22'b0000000101010001111011,
    22'b0000000110011001100110,
    22'b0000000111001100110011,
    22'b0000001000000000000000,
    22'b0000001000011110101110,
    22'b0000001000101000111101,
    22'b0000001000011110101110,
    22'b0000001000000000000000,
    22'b0000000111010111000011,
    22'b0000000110100011110110,
    22'b0000000101100110011010,
    22'b0000000100001010001111,
    22'b0000000011001100110011,
    22'b0000000010000101001000,
    22'b0000000001000111101100,
    22'b0000000000000000000000,
    22'b0000000001010001111011,
    22'b0000000001011100001010,
    22'b0000000001110000101001,
    22'b0000000010011001100110,
    22'b0000000010101110000101,
    22'b0000000011001100110011,
    22'b0000000011101011100001,
    22'b0000000100001010001111,
    22'b0000000100011110101110,
    22'b0000000100101000111101,
    22'b0000000101000111101100,
    22'b0000000101110000101001,
    22'b0000000101111010111000,
    22'b0000000101100110011010,
    22'b0000000100111101011100,
    22'b0000000100011110101110,
    22'b0000000101011100001010,
    22'b0000000111001100110011,
    22'b0000001010100011110110,
    22'b0000001100101000111101,
    22'b0000001110001111010111,
    22'b0000001111000010100100,
    22'b0000001111010111000011,
    22'b0000001111010111000011,
    22'b0000001111100001010010,
    22'b0000010000001010001111,
    22'b0000010001010001111011,
    22'b0000010011001100110011,
    22'b0000010100101000111101,
    22'b0000010110000101001000,
    22'b0000010111010111000011,
    22'b0000011001010001111011,
    22'b0000011010111000010100,
    22'b0000011100010100011111,
    22'b0000011100101000111101,
    22'b0000011100110011001101,
    22'b0000100000000000000000,
    22'b0000100010001111010111,
    22'b0000100011100001010010,
    22'b0000100100011110101110,
    22'b0000100101110000101001,
    22'b0000100110100011110110,
    22'b0000100111100001010010,
    22'b0000101000110011001101,
    22'b0000101010100011110110,
    22'b0000101101010001111011,
    22'b0000101111000010100100,
    22'b0000110001010001111011,
    22'b0000110100110011001101,
    22'b0000111000101000111101,
    22'b0000111100111101011100,
    22'b0001000000101000111101,
    22'b0001000100011110101110,
    22'b0001001010111000010100,
    22'b0001001111100001010010,
    22'b0001010010001111010111,
    22'b0001010010011001100110,
    22'b0001010000001010001111,
    22'b0001001010100011110110,
    22'b0001000101010001111011,
    22'b0000111111110101110001,
    22'b0000111010100011110110,
    22'b0000110100110011001101,
    22'b0000110001110000101001,
    22'b0000101111110101110001,
    22'b0000101110011001100110,
    22'b0000101100011110101110,
    22'b0000101001110000101001,
    22'b0000100111001100110011,
    22'b0000100100011110101110,
    22'b0000011111101011100001,
    22'b0000011100000000000000,
    22'b0000011000110011001101,
    22'b0000010110011001100110,
    22'b0000010100111101011100,
    22'b0000010011110101110001,
    22'b0000010011110101110001,
    22'b0000010100101000111101,
    22'b0000010101111010111000,
    22'b0000011000111101011100,
    22'b0000011011101011100001,
    22'b0000011110101110000101,
    22'b0000100001010001111011,
    22'b0000100011001100110011,
    22'b0000100100110011001101,
    22'b0000100101010001111011,
    22'b0000100100111101011100,
    22'b0000100100000000000000,
    22'b0000100001100110011010,
    22'b0000011111100001010010,
    22'b0000011101010001111011,
    22'b0000011011000010100100,
    22'b0000011000110011001101,
    22'b0000010110101110000101,
    22'b0000010101111010111000,
    22'b0000010101110000101001,
    22'b0000010110001111010111,
    22'b0000010110101110000101,
    22'b0000010111001100110011,
    22'b0000010111001100110011,
    22'b0000010110100011110110,
    22'b0000010101110000101001,
    22'b0000010101000111101100,
    22'b0000010011110101110001,
    22'b0000010001110000101001,
    22'b0000001111010111000011,
    22'b0000001100110011001101,
    22'b0000001010101110000101,
    22'b0000001000011110101110,
    22'b0000000111010111000011,
    22'b0000000110011001100110,
    22'b0000000101110000101001,
    22'b0000000100111101011100,
    22'b0000000100010100011111,
    22'b0000000011001100110011,
    22'b0000000001100110011010,
    22'b1111111111101011100001,
    22'b1111111100111101011100,
    22'b1111111010101110000101,
    22'b1111111000101000111101,
    22'b1111110111000010100100,
    22'b1111110110100011110110,
    22'b1111110101000111101100,
    22'b1111110100011110101110,
    22'b1111110110000101001000,
    22'b1111111000001010001111,
    22'b1111111000001010001111,
    22'b1111110100111101011100,
    22'b1111110011010111000011,
    22'b1111110010011001100110,
    22'b1111110001011100001010,
    22'b1111101111110101110001,
    22'b1111101111000010100100,
    22'b1111101101011100001010,
    22'b1111101010111000010100,
    22'b1111100111110101110001,
    22'b1111100011101011100001,
    22'b1111100000011110101110,
    22'b1111011101010001111011,
    22'b1111011010111000010100,
    22'b1111011001000111101100,
    22'b1111010111100001010010,
    22'b1111010111000010100100,
    22'b1111010110111000010100,
    22'b1111010111100001010010,
    22'b1111011000001010001111,
    22'b1111011000101000111101,
    22'b1111011000110011001101,
    22'b1111011000011110101110,
    22'b1111010111110101110001,
    22'b1111010110000101001000,
    22'b1111010100111101011100,
    22'b1111010100000000000000,
    22'b1111010011100001010010,
    22'b1111010011101011100001,
    22'b1111010100101000111101,
    22'b1111010101111010111000,
    22'b1111010111010111000011,
    22'b1111011000011110101110,
    22'b1111011001011100001010,
    22'b1111011001011100001010,
    22'b1111011000111101011100,
    22'b1111011000001010001111,
    22'b1111010110100011110110,
    22'b1111010101011100001010,
    22'b1111010100010100011111,
    22'b1111010100011110101110,
    22'b1111010110000101001000,
    22'b1111011001110000101001,
    22'b1111011110111000010100,
    22'b1111100011010111000011,
    22'b1111101000000000000000,
    22'b1111101100111101011100,
    22'b1111101110101110000101,
    22'b1111101111010111000011,
    22'b1111101111101011100001,
    22'b1111110000000000000000,
    22'b1111110000011110101110,
    22'b1111110000111101011100,
    22'b1111110001010001111011,
    22'b1111110001011100001010,
    22'b1111110001010001111011,
    22'b1111110000101000111101,
    22'b1111101111101011100001,
    22'b1111101110000101001000,
    22'b1111101100110011001101,
    22'b1111101011100001010010,
    22'b1111101010100011110110,
    22'b1111101010000101001000,
    22'b1111101011100001010010,
    22'b1111101110001111010111,
    22'b1111101111010111000011,
    22'b1111101111010111000011,
    22'b1111110000010100011111,
    22'b1111110000111101011100,
    22'b1111110010001111010111,
    22'b1111110011101011100001,
    22'b1111110100110011001101,
    22'b1111110100010100011111,
    22'b1111110011110101110001,
    22'b1111110001110000101001,
    22'b1111101111100001010010,
    22'b1111101101111010111000,
    22'b1111101100010100011111,
    22'b1111101001111010111000,
    22'b1111101000011110101110,
    22'b1111100111000010100100,
    22'b1111100101111010111000,
    22'b1111100101000111101100,
    22'b1111100100111101011100,
    22'b1111100101011100001010,
    22'b1111100111101011100001,
    22'b1111101100010100011111,
    22'b1111110000101000111101,
    22'b1111110101000111101100,
    22'b1111111000011110101110,
    22'b1111111010000101001000,
    22'b1111111001010001111011,
    22'b1111110111010111000011,
    22'b1111110101111010111000,
    22'b1111110010100011110110,
    22'b1111110000010100011111,
    22'b1111101100111101011100,
    22'b1111101001011100001010,
    22'b1111101001110000101001,
    22'b1111101101000111101100,
    22'b1111110000101000111101,
    22'b1111110011000010100100,
    22'b1111110100101000111101,
    22'b1111110101000111101100,
    22'b1111110100110011001101,
    22'b1111110011101011100001,
    22'b1111110001010001111011,
    22'b1111101111010111000011,
    22'b1111101110011001100110,
    22'b1111101110000101001000,
    22'b1111101110001111010111,
    22'b1111101110100011110110,
    22'b1111101110001111010111,
    22'b1111101000001010001111,
    22'b1111100111100001010010,
    22'b1111100111010111000011,
    22'b1111100111100001010010,
    22'b1111101000001010001111,
    22'b1111101000110011001101,
    22'b1111101001000111101100,
    22'b1111101001011100001010,
    22'b1111101001010001111011,
    22'b1111101001000111101100,
    22'b1111101000110011001101,
    22'b1111101000101000111101,
    22'b1111101000101000111101,
    22'b1111101000101000111101,
    22'b1111101000011110101110,
    22'b1111101000101000111101,
    22'b1111101000101000111101,
    22'b1111101000111101011100,
    22'b1111101001010001111011,
    22'b1111101001110000101001,
    22'b1111101010001111010111,
    22'b1111101010111000010100,
    22'b1111101011101011100001,
    22'b1111101101000111101100,
    22'b1111101110011001100110,
    22'b1111110000101000111101,
    22'b1111110100110011001101,
    22'b1111111001110000101001,
    22'b1111111101000111101100,
    22'b1111111110100011110110,
    22'b1111111111101011100001,
    22'b1111111101100110011010,
    22'b1111111011010111000011,
    22'b1111111001110000101001,
    22'b1111111000011110101110,
    22'b1111110111100001010010,
    22'b1111110110011001100110,
    22'b1111110100010100011111,
    22'b1111110000110011001101,
    22'b1111101101111010111000,
    22'b1111101001111010111000,
    22'b1111100101011100001010,
    22'b1111011111101011100001,
    22'b1111011100001010001111,
    22'b1111011001110000101001,
    22'b1111011000010100011111,
    22'b1111010111000010100100,
    22'b1111010110111000010100,
    22'b1111010110111000010100,
    22'b1111010111010111000011,
    22'b1111011000010100011111,
    22'b1111011000111101011100,
    22'b1111011000111101011100,
    22'b1111011000011110101110,
    22'b1111010111110101110001,
    22'b1111010111100001010010,
    22'b1111010111101011100001,
    22'b1111011000011110101110,
    22'b1111011001011100001010,
    22'b1111011010100011110110,
    22'b1111011011110101110001,
    22'b1111011101000111101100,
    22'b1111011110100011110110,
    22'b1111100000001010001111,
    22'b1111100001110000101001,
    22'b1111100011110101110001,
    22'b1111101000011110101110,
    22'b1111101001000111101100,
    22'b1111101001111010111000,
    22'b1111101010100011110110,
    22'b1111101011000010100100,
    22'b1111101011010111000011,
    22'b1111101011000010100100,
    22'b1111101010001111010111,
    22'b1111101000111101011100,
    22'b1111100111101011100001,
    22'b1111100110001111010111,
    22'b1111100101011100001010,
    22'b1111100101000111101100,
    22'b1111100100110011001101,
    22'b1111100100101000111101,
    22'b1111100100101000111101,
    22'b1111100100111101011100,
    22'b1111100110001111010111,
    22'b1111100111100001010010,
    22'b1111101001010001111011,
    22'b1111101011000010100100,
    22'b1111101100011110101110,
    22'b1111101101111010111000,
    22'b1111101110111000010100,
    22'b1111110000000000000000,
    22'b1111110001010001111011,
    22'b1111110011001100110011,
    22'b1111110100111101011100,
    22'b1111110110100011110110,
    22'b1111110111110101110001,
    22'b1111111000111101011100,
    22'b1111111001100110011010,
    22'b1111111010000101001000,
    22'b1111111010111000010100,
    22'b1111111100000000000000,
    22'b1111111100011110101110,
    22'b1111111100111101011100,
    22'b1111111101010001111011,
    22'b1111111100111101011100,
    22'b1111111100011110101110,
    22'b1111111100000000000000,
    22'b1111111011110101110001,
    22'b1111111011110101110001,
    22'b1111111011101011100001,
    22'b1111111011101011100001,
    22'b1111111011100001010010,
    22'b1111111011001100110011,
    22'b1111111011001100110011,
    22'b1111111011001100110011,
    22'b1111111011101011100001,
    22'b1111111100000000000000,
    22'b1111111100011110101110,
    22'b1111111100111101011100,
    22'b1111111111101011100001,
    22'b0000000000001010001111,
    22'b0000000000011110101110,
    22'b0000000000110011001101,
    22'b0000000001010001111011,
    22'b0000000001011100001010,
    22'b0000000001100110011010,
    22'b0000000001111010111000,
    22'b0000000010001111010111,
    22'b0000000010111000010100,
    22'b0000000011100001010010,
    22'b0000000100000000000000,
    22'b0000000100011110101110,
    22'b0000000101000111101100,
    22'b0000000101100110011010,
    22'b0000000110000101001000,
    22'b0000000110100011110110,
    22'b0000000111000010100100,
    22'b0000000111100001010010,
    22'b0000000111110101110001,
    22'b0000000111101011100001,
    22'b0000000111100001010010,
    22'b0000000111110101110001,
    22'b0000001000001010001111,
    22'b0000001000001010001111,
    22'b0000001000001010001111,
    22'b0000001000000000000000,
    22'b0000000111010111000011,
    22'b0000000110001111010111,
    22'b0000000100110011001101,
    22'b0000000011001100110011,
    22'b0000000000110011001101,
    22'b1111111110101110000101,
    22'b1111111100101000111101,
    22'b1111111011000010100100,
    22'b1111111001000111101100,
    22'b1111110111101011100001,
    22'b1111110110011001100110,
    22'b1111110101010001111011,
    22'b1111110010101110000101,
    22'b1111110000111101011100,
    22'b1111101111101011100001,
    22'b1111101110011001100110,
    22'b1111101100101000111101,
    22'b1111101011001100110011,
    22'b1111101001100110011010,
    22'b1111101000000000000000,
    22'b1111100111001100110011,
    22'b1111100110001111010111,
    22'b1111100101100110011010,
    22'b1111100101010001111011,
    22'b1111100101100110011010,
    22'b1111100101000111101100,
    22'b1111100110101110000101,
    22'b1111101001000111101100,
    22'b1111101100010100011111,
    22'b1111110000111101011100,
    22'b1111110111001100110011,
    22'b0000000010000101001000,
    22'b0000010011100001010010,
    22'b0000011111000010100100,
    22'b0000100101010001111011,
    22'b0000100111001100110011,
    22'b0000100111100001010010,
    22'b0000100101111010111000,
    22'b0000100101100110011010,
    22'b0000100100110011001101,
    22'b0000100010000101001000,
    22'b0000011101100110011010,
    22'b0000010110000101001000,
    22'b0000010000111101011100,
    22'b0000001101111010111000,
    22'b0000001001111010111000,
    22'b0000001000010100011111,
    22'b0000001000001010001111,
    22'b0000001000000000000000,
    22'b0000000111100001010010,
    22'b0000000110101110000101,
    22'b0000000101011100001010,
    22'b0000000100110011001101,
    22'b0000000100101000111101,
    22'b0000000100011110101110,
    22'b0000000100110011001101,
    22'b0000000110011001100110,
    22'b0000001011110101110001,
    22'b0000010100000000000000,
    22'b0000011011101011100001,
    22'b0000011111100001010010,
    22'b0000011001111010111000,
    22'b0000010011001100110011,
    22'b0000001100111101011100,
    22'b0000000111101011100001,
    22'b0000000001110000101001,
    22'b1111111110101110000101,
    22'b1111111100011110101110,
    22'b1111111010000101001000,
    22'b1111110101011100001010,
    22'b1111110001000111101100,
    22'b1111101100110011001101,
    22'b1111101010101110000101,
    22'b1111101011010111000011,
    22'b1111101011010111000011,
    22'b1111101011001100110011,
    22'b1111101011001100110011,
    22'b1111101010111000010100,
    22'b1111101010001111010111,
    22'b1111101000111101011100,
    22'b1111100110100011110110,
    22'b1111100100110011001101,
    22'b1111100001111010111000,
    22'b1111011111100001010010,
    22'b1111011110001111010111,
    22'b1111011111010111000011,
    22'b1111100001000111101100,
    22'b1111100010101110000101,
    22'b1111100011101011100001,
    22'b1111100100101000111101,
    22'b1111100100110011001101,
    22'b1111100100011110101110,
    22'b1111100011101011100001,
    22'b1111100010111000010100,
    22'b1111100001100110011010,
    22'b1111011111001100110011,
    22'b1111011100101000111101,
    22'b1111011001111010111000,
    22'b1111010111110101110001,
    22'b1111010110001111010111,
    22'b1111011000111101011100,
    22'b1111011110101110000101,
    22'b1111011111000010100100,
    22'b1111011111100001010010,
    22'b1111011111110101110001,
    22'b1111011010000101001000,
    22'b1111010111110101110001,
    22'b1111010101110000101001,
    22'b1111010011001100110011,
    22'b1111010001011100001010,
    22'b1111010000000000000000,
    22'b1111001110011001100110,
    22'b1111001101100110011010,
    22'b1111001101010001111011,
    22'b1111001101000111101100,
    22'b1111001100111101011100,
    22'b1111001100110011001101,
    22'b1111001100010100011111,
    22'b1111001100000000000000,
    22'b1111001011010111000011,
    22'b1111001011000010100100,
    22'b1111001010111000010100,
    22'b1111001010111000010100,
    22'b1111001011010111000011,
    22'b1111001011110101110001,
    22'b1111001100101000111101,
    22'b1111001101010001111011,
    22'b1111001110011001100110,
    22'b1111001111010111000011,
    22'b1111010000010100011111,
    22'b1111010001011100001010,
    22'b1111010010101110000101,
    22'b1111010011100001010010,
    22'b1111010100010100011111,
    22'b1111010101000111101100,
    22'b1111010110011001100110,
    22'b1111010111100001010010,
    22'b1111011000001010001111,
    22'b1111011000011110101110,
    22'b1111011000010100011111,
    22'b1111011000011110101110,
    22'b1111011000110011001101,
    22'b1111011001000111101100,
    22'b1111011001011100001010,
    22'b1111011001010001111011,
    22'b1111011001000111101100,
    22'b1111011000111101011100,
    22'b1111011000011110101110,
    22'b1111011000010100011111,
    22'b1111011000001010001111,
    22'b1111011000010100011111,
    22'b1111011000101000111101,
    22'b1111011000111101011100,
    22'b1111011001000111101100,
    22'b1111011001111010111000,
    22'b1111011011000010100100,
    22'b1111011100000000000000,
    22'b1111011100011110101110,
    22'b1111011101010001111011,
    22'b1111011101110000101001,
    22'b1111011110001111010111,
    22'b1111011110100011110110,
    22'b1111011111001100110011,
    22'b1111100000000000000000,
    22'b1111100001010001111011,
    22'b1111100011101011100001,
    22'b1111100110001111010111,
    22'b1111101000110011001101,
    22'b1111101011010111000011,
    22'b1111111010000101001000,
    22'b1111111110011001100110,
    22'b0000000001010001111011,
    22'b0000000010100011110110,
    22'b0000000110101110000101,
    22'b0000001011010111000011,
    22'b0000001110111000010100,
    22'b0000010000110011001101,
    22'b0000010001111010111000,
    22'b0000010001100110011010,
    22'b0000010000111101011100,
    22'b0000010001011100001010,
    22'b0000010001000111101100,
    22'b0000001111000010100100,
    22'b0000001001100110011010,
    22'b0000000010101110000101,
    22'b1111111110111000010100,
    22'b1111111101110000101001,
    22'b1111111110011001100110,
    22'b0000000000011110101110,
    22'b0000000011001100110011,
    22'b0000000110001111010111,
    22'b0000001011110101110001,
    22'b0000010000000000000000,
    22'b0000010011101011100001,
    22'b0000010111000010100100,
    22'b0000011010000101001000,
    22'b0000011101111010111000,
    22'b0000100000111101011100,
    22'b0000100011101011100001,
    22'b0000100101100110011010,
    22'b0000100110111000010100,
    22'b0000101000110011001101,
    22'b0000101010001111010111,
    22'b0000101010001111010111,
    22'b0000101001000111101100,
    22'b0000100111101011100001,
    22'b0000100111100001010010,
    22'b0000100111000010100100,
    22'b0000100101110000101001,
    22'b0000100100001010001111,
    22'b0000100010001111010111,
    22'b0000100010100011110110,
    22'b0000100001111010111000,
    22'b0000100001000111101100,
    22'b0000100000001010001111,
    22'b0000011110101110000101,
    22'b0000011110011001100110,
    22'b0000011100011110101110,
    22'b0000011010000101001000,
    22'b0000010111001100110011,
    22'b0000010011001100110011,
    22'b0000010000101000111101,
    22'b0000001110101110000101,
    22'b0000001101100110011010,
    22'b0000001100011110101110,
    22'b0000001101110000101001,
    22'b0000001111000010100100,
    22'b0000010000110011001101,
    22'b0000010010011001100110,
    22'b0000010100101000111101,
    22'b0000010110101110000101,
    22'b0000010111110101110001,
    22'b0000010111110101110001,
    22'b0000010111100001010010,
    22'b0000010111000010100100,
    22'b0000010110111000010100,
    22'b0000010110101110000101,
    22'b0000010111100001010010,
    22'b0000011001111010111000,
    22'b0000011001010001111011,
    22'b0000010111100001010010,
    22'b0000010111000010100100,
    22'b0000010100111101011100,
    22'b0000010001111010111000,
    22'b0000010000000000000000,
    22'b0000001111101011100001,
    22'b0000001111100001010010,
    22'b0000010001100110011010,
    22'b0000010000010100011111,
    22'b0000010010001111010111,
    22'b0000010100110011001101,
    22'b0000010110011001100110,
    22'b0000011000010100011111,
    22'b0000010100001010001111,
    22'b0000010000011110101110,
    22'b0000001101010001111011,
    22'b0000001010011001100110,
    22'b0000001111010111000011,
    22'b0000010101000111101100,
    22'b0000010011110101110001,
    22'b0000010000101000111101,
    22'b0000001110111000010100,
    22'b0000001100111101011100,
    22'b0000001001010001111011,
    22'b0000000101111010111000,
    22'b0000000100001010001111,
    22'b0000000100101000111101,
    22'b0000000101111010111000,
    22'b0000000111001100110011,
    22'b0000001000010100011111,
    22'b0000001000111101011100,
    22'b0000001000111101011100,
    22'b0000001000011110101110,
    22'b0000001000001010001111,
    22'b0000001000000000000000,
    22'b0000000111110101110001,
    22'b0000000111101011100001,
    22'b0000000111100001010010,
    22'b0000000111101011100001,
    22'b0000001000010100011111,
    22'b0000001001110000101001,
    22'b0000001010100011110110,
    22'b0000001011000010100100,
    22'b0000001011001100110011,
    22'b0000001011100001010010,
    22'b0000001101100110011010,
    22'b0000001110101110000101,
    22'b0000010000000000000000,
    22'b0000010000111101011100,
    22'b0000010001100110011010,
    22'b0000010001111010111000,
    22'b0000010001100110011010,
    22'b0000010001010001111011,
    22'b0000010000111101011100,
    22'b0000010000110011001101,
    22'b0000010000010100011111,
    22'b0000001111101011100001,
    22'b0000001111000010100100,
    22'b0000001101111010111000,
    22'b0000001100111101011100,
    22'b0000001011100001010010,
    22'b0000001010111000010100,
    22'b0000001010100011110110,
    22'b0000001010100011110110,
    22'b0000001010001111010111,
    22'b0000001001111010111000,
    22'b0000001001111010111000,
    22'b0000001001111010111000,
    22'b0000001010001111010111,
    22'b0000001011000010100100,
    22'b0000001011100001010010,
    22'b0000001011101011100001,
    22'b0000001011010111000011,
    22'b0000001011001100110011,
    22'b0000001010100011110110,
    22'b0000001001011100001010,
    22'b0000001000011110101110,
    22'b0000000111100001010010,
    22'b0000000110100011110110,
    22'b0000000101100110011010,
    22'b0000000100101000111101,
    22'b0000000100010100011111,
    22'b0000000100110011001101,
    22'b0000000101011100001010,
    22'b0000000110101110000101,
    22'b0000001001110000101001,
    22'b0000001100000000000000,
    22'b0000001110001111010111,
    22'b0000001110111000010100,
    22'b0000010000000000000000,
    22'b0000010001010001111011,
    22'b0000010000111101011100,
    22'b0000010000111101011100,
    22'b0000010001011100001010,
    22'b0000010010001111010111,
    22'b0000010011000010100100,
    22'b0000010011101011100001,
    22'b0000010100010100011111,
    22'b0000010100111101011100,
    22'b0000010101111010111000,
    22'b0000010110011001100110,
    22'b0000010101111010111000,
    22'b0000010100101000111101,
    22'b0000010101010001111011,
    22'b0000010101000111101100,
    22'b0000010011101011100001,
    22'b0000010010011001100110,
    22'b0000010010000101001000,
    22'b0000010001111010111000,
    22'b0000010010000101001000,
    22'b0000010010111000010100,
    22'b0000010100000000000000,
    22'b0000010100110011001101,
    22'b0000010100101000111101,
    22'b0000010100011110101110,
    22'b0000010100000000000000,
    22'b0000010011001100110011,
    22'b0000010010000101001000,
    22'b0000010000011110101110,
    22'b0000001111110101110001,
    22'b0000001111101011100001,
    22'b0000010000000000000000,
    22'b0000010000010100011111,
    22'b0000010000101000111101,
    22'b0000010000010100011111,
    22'b0000001111101011100001,
    22'b0000001110100011110110,
    22'b0000001100110011001101,
    22'b0000001011100001010010,
    22'b0000001010011001100110,
    22'b0000001001100110011010,
    22'b0000001000110011001101,
    22'b0000001000010100011111,
    22'b0000001000011110101110,
    22'b0000001001000111101100,
    22'b0000001001011100001010,
    22'b0000001010111000010100,
    22'b0000001101011100001010,
    22'b0000010000000000000000,
    22'b0000010010111000010100,
    22'b0000010100101000111101,
    22'b0000010110011001100110,
    22'b0000010111001100110011,
    22'b0000011000101000111101,
    22'b0000011000110011001101,
    22'b0000011000001010001111,
    22'b0000010111000010100100,
    22'b0000010110000101001000,
    22'b0000010100110011001101,
    22'b0000010011110101110001,
    22'b0000010011000010100100,
    22'b0000010001011100001010,
    22'b0000010000101000111101,
    22'b0000010000001010001111,
    22'b0000001111110101110001,
    22'b0000001111101011100001,
    22'b0000001111010111000011,
    22'b0000001111000010100100,
    22'b0000001110011001100110,
    22'b0000001101110000101001,
    22'b0000001100101000111101,
    22'b0000001010100011110110,
    22'b0000001000001010001111,
    22'b0000000101111010111000,
    22'b0000000100000000000000,
    22'b0000000010001111010111,
    22'b1111111111110101110001,
    22'b1111111110100011110110,
    22'b1111111101000111101100,
    22'b1111111100010100011111,
    22'b1111111011010111000011,
    22'b1111111011000010100100,
    22'b1111111000011110101110,
    22'b1111110101010001111011,
    22'b1111110001011100001010,
    22'b1111101101010001111011,
    22'b1111101101011100001010,
    22'b1111110000000000000000,
    22'b1111110011101011100001,
    22'b1111111010111000010100,
    22'b0000000000000000000000,
    22'b0000000110001111010111,
    22'b0000001100111101011100,
    22'b0000010010000101001000,
    22'b0000010100111101011100,
    22'b0000010101010001111011,
    22'b0000010100000000000000,
    22'b0000010001100110011010,
    22'b0000001110111000010100,
    22'b0000001011100001010010,
    22'b0000001001000111101100,
    22'b0000000111000010100100,
    22'b0000000100110011001101,
    22'b0000000000111101011100,
    22'b1111111100010100011111,
    22'b1111110111110101110001,
    22'b1111110100001010001111,
    22'b1111110001110000101001,
    22'b1111110000101000111101,
    22'b1111110010111000010100,
    22'b1111110101111010111000,
    22'b1111111000010100011111,
    22'b1111111010011001100110,
    22'b1111111010111000010100,
    22'b1111111011001100110011,
    22'b1111111011101011100001,
    22'b1111111100011110101110,
    22'b1111111111001100110011,
    22'b0000000001011100001010,
    22'b0000000011010111000011,
    22'b0000000101000111101100,
    22'b0000000110011001100110,
    22'b0000000110101110000101,
    22'b0000000111000010100100,
    22'b0000000111100001010010,
    22'b0000001000011110101110,
    22'b0000001001010001111011,
    22'b0000001010011001100110,
    22'b0000001011100001010010,
    22'b0000001100110011001101,
    22'b0000001110111000010100,
    22'b0000010000101000111101,
    22'b0000010010011001100110,
    22'b0000010100010100011111,
    22'b0000010110100011110110,
    22'b0000010111110101110001,
    22'b0000011000101000111101,
    22'b0000011001011100001010,
    22'b0000011010000101001000,
    22'b0000011010100011110110,
    22'b0000011010111000010100,
    22'b0000011010001111010111,
    22'b0000011011001100110011,
    22'b0000011011101011100001,
    22'b0000011100010100011111,
    22'b0000011100111101011100,
    22'b0000011101110000101001,
    22'b0000011110111000010100,
    22'b0000100000110011001101,
    22'b0000100001110000101001,
    22'b0000100010001111010111,
    22'b0000100100001010001111,
    22'b0000100101100110011010,
    22'b0000101000101000111101,
    22'b0000101100001010001111,
    22'b0000110001100110011010,
    22'b0000110111000010100100,
    22'b0000111101100110011010,
    22'b0001000001100110011010,
    22'b0001000001111010111000,
    22'b0000111000000000000000,
    22'b0000011101100110011010,
    22'b0000001101110000101001,
    22'b0000001011000010100100,
    22'b0000010100101000111101,
    22'b0000011100000000000000,
    22'b0000011100110011001101,
    22'b0000011000110011001101,
    22'b0000010111100001010010,
    22'b0000011100001010001111,
    22'b0000100010101110000101,
    22'b0000101000101000111101,
    22'b0000101100101000111101,
    22'b0000101101011100001010,
    22'b0000101001011100001010,
    22'b0000100100101000111101,
    22'b0000011111101011100001,
    22'b0000011100000000000000,
    22'b0000011001011100001010,
    22'b0000011000111101011100,
    22'b0000011001011100001010,
    22'b0000011010011001100110,
    22'b0000011011100001010010,
    22'b0000011100111101011100,
    22'b0000011101011100001010,
    22'b0000011101100110011010,
    22'b0000011101011100001010,
    22'b0000011100011110101110,
    22'b0000011011010111000011,
    22'b0000011010000101001000,
    22'b0000011001000111101100,
    22'b0000011000010100011111,
    22'b0000010111100001010010,
    22'b0000010110001111010111,
    22'b0000010101000111101100,
    22'b0000010011000010100100,
    22'b0000010001100110011010,
    22'b0000010000010100011111,
    22'b0000001111101011100001,
    22'b0000001110101110000101,
    22'b0000001110000101001000,
    22'b0000001101100110011010,
    22'b0000001101010001111011,
    22'b0000001100101000111101,
    22'b0000001011010111000011,
    22'b0000001010000101001000,
    22'b0000001000110011001101,
    22'b0000000111101011100001,
    22'b0000000111000010100100,
    22'b0000000110111000010100,
    22'b0000000111010111000011,
    22'b0000000111110101110001,
    22'b0000001000011110101110,
    22'b0000001000111101011100,
    22'b0000001001110000101001,
    22'b0000001010011001100110,
    22'b0000001010111000010100,
    22'b0000001011000010100100,
    22'b0000001010101110000101,
    22'b0000001010011001100110,
    22'b0000001001111010111000,
    22'b0000001001010001111011,
    22'b0000001000101000111101,
    22'b0000001000001010001111,
    22'b0000000111110101110001,
    22'b0000000111100001010010,
    22'b0000000111010111000011,
    22'b0000000111001100110011,
    22'b0000000110111000010100,
    22'b0000000101111010111000,
    22'b0000000100010100011111,
    22'b0000000010101110000101,
    22'b0000000001010001111011,
    22'b1111111111110101110001,
    22'b1111111110100011110110,
    22'b1111111100110011001101,
    22'b1111111011101011100001,
    22'b1111111010100011110110,
    22'b1111111001011100001010,
    22'b1111110111110101110001,
    22'b1111110110100011110110,
    22'b1111110101010001111011,
    22'b1111110100001010001111,
    22'b1111110010101110000101,
    22'b1111110001110000101001,
    22'b1111110000111101011100,
    22'b1111110000001010001111,
    22'b1111101111101011100001,
    22'b1111101111001100110011,
    22'b1111101110111000010100,
    22'b1111101110101110000101,
    22'b1111101110101110000101,
    22'b1111101110101110000101,
    22'b1111101110101110000101,
    22'b1111101110100011110110,
    22'b1111101110011001100110,
    22'b1111101110001111010111,
    22'b1111101110000101001000,
    22'b1111101101111010111000,
    22'b1111101101011100001010,
    22'b1111101101000111101100,
    22'b1111101100101000111101,
    22'b1111101100110011001101,
    22'b1111101101000111101100,
    22'b1111101101111010111000,
    22'b1111101111100001010010,
    22'b1111110000011110101110,
    22'b1111110001010001111011,
    22'b1111110001110000101001,
    22'b1111110001010001111011,
    22'b1111110000001010001111,
    22'b1111101110101110000101,
    22'b1111101101010001111011,
    22'b1111101011101011100001,
    22'b1111101010111000010100,
    22'b1111101010100011110110,
    22'b1111101010011001100110,
    22'b1111101010100011110110,
    22'b1111101011001100110011,
    22'b1111101100000000000000,
    22'b1111101100110011001101,
    22'b1111101101110000101001,
    22'b1111101110111000010100,
    22'b1111101111101011100001,
    22'b1111110000001010001111,
    22'b1111110000011110101110,
    22'b1111110000111101011100,
    22'b1111110001010001111011,
    22'b1111110001110000101001,
    22'b1111110010011001100110,
    22'b1111110011101011100001,
    22'b1111110100101000111101,
    22'b1111110101100110011010,
    22'b1111110110011001100110,
    22'b1111110111010111000011,
    22'b1111110111110101110001,
    22'b1111110111110101110001,
    22'b1111110111101011100001,
    22'b1111110111001100110011,
    22'b1111110110111000010100,
    22'b1111110110100011110110,
    22'b1111110110011001100110,
    22'b1111110110100011110110,
    22'b1111110110111000010100,
    22'b1111110111100001010010,
    22'b1111111000101000111101,
    22'b1111111010100011110110,
    22'b1111111100010100011111,
    22'b1111111101111010111000,
    22'b1111111111000010100100,
    22'b1111111111110101110001,
    22'b0000000000000000000000,
    22'b1111111111101011100001,
    22'b1111111111100001010010,
    22'b1111111111010111000011,
    22'b1111111111010111000011,
    22'b1111111111101011100001,
    22'b1111111111101011100001,
    22'b1111111111000010100100,
    22'b1111111110001111010111,
    22'b1111111011101011100001,
    22'b1111110111110101110001,
    22'b1111110010101110000101,
    22'b1111101110011001100110,
    22'b1111101010011001100110,
    22'b1111100111000010100100,
    22'b1111100011100001010010,
    22'b1111100001100110011010,
    22'b1111100000010100011111,
    22'b1111011111010111000011,
    22'b1111011110101110000101,
    22'b1111011110011001100110,
    22'b1111011110100011110110,
    22'b1111011111001100110011,
    22'b1111100000000000000000,
    22'b1111100000111101011100,
    22'b1111100010000101001000,
    22'b1111100011001100110011,
    22'b1111100100110011001101,
    22'b1111100101110000101001,
    22'b1111100110101110000101,
    22'b1111100111100001010010,
    22'b1111101000110011001101,
    22'b1111101010000101001000,
    22'b1111101011100001010010,
    22'b1111101101010001111011,
    22'b1111101111100001010010,
    22'b1111110000111101011100,
    22'b1111110001000111101100,
    22'b1111110000001010001111,
    22'b1111101101011100001010,
    22'b1111101011000010100100,
    22'b1111101000001010001111,
    22'b1111100101000111101100,
    22'b1111011111101011100001,
    22'b1111011010101110000101,
    22'b1111010101111010111000,
    22'b1111010001010001111011,
    22'b1111001011100001010010,
    22'b1111000111101011100001,
    22'b1111000100101000111101,
    22'b1111000001110000101001,
    22'b1111000011000010100100,
    22'b1111000101000111101100,
    22'b1111000111100001010010,
    22'b1111001001011100001010,
    22'b1111001011110101110001,
    22'b1111001110101110000101,
    22'b1111010010000101001000,
    22'b1111010100101000111101,
    22'b1111010110101110000101,
    22'b1111011000011110101110,
    22'b1111011010011001100110,
    22'b1111011011101011100001,
    22'b1111011101000111101100,
    22'b1111011110100011110110,
    22'b1111100000011110101110,
    22'b1111100001011100001010,
    22'b1111100010011001100110,
    22'b1111100011001100110011,
    22'b1111100100001010001111,
    22'b1111100100111101011100,
    22'b1111100101110000101001,
    22'b1111100110011001100110,
    22'b1111100111010111000011,
    22'b1111100111110101110001,
    22'b1111101000011110101110,
    22'b1111101000111101011100,
    22'b1111101001000111101100,
    22'b1111101001000111101100,
    22'b1111101000111101011100,
    22'b1111101000101000111101,
    22'b1111101000010100011111,
    22'b1111100111110101110001,
    22'b1111100111100001010010,
    22'b1111100111000010100100,
    22'b1111101000000000000000,
    22'b1111101010000101001000,
    22'b1111101011101011100001,
    22'b1111101011010111000011,
    22'b1111100110101110000101,
    22'b1111011111110101110001,
    22'b1111011000000000000000,
    22'b1111001101000111101100,
    22'b1111000100001010001111,
    22'b1110111011001100110011,
    22'b1110110000001010001111,
    22'b1110101001100110011010,
    22'b1110100101000111101100,
    22'b1110100011000010100100,
    22'b1110100100000000000000,
    22'b1110100111000010100100,
    22'b1110101010011001100110,
    22'b1110101110000101001000,
    22'b1110110011010111000011,
    22'b1110110111010111000011,
    22'b1110111100000000000000,
    22'b1111000000111101011100,
    22'b1111000111100001010010,
    22'b1111010111000010100100,
    22'b1111011010000101001000,
    22'b1111011101111010111000,
    22'b1111100000011110101110,
    22'b1111100010101110000101,
    22'b1111100100011110101110,
    22'b1111100110000101001000,
    22'b1111100111000010100100,
    22'b1111100111110101110001,
    22'b1111101000110011001101,
    22'b1111101001100110011010,
    22'b1111101010011001100110,
    22'b1111101011001100110011,
    22'b1111101100011110101110,
    22'b1111101101011100001010,
    22'b1111101110101110000101,
    22'b1111110000001010001111,
    22'b1111110010000101001000,
    22'b1111110011101011100001,
    22'b1111110101011100001010,
    22'b1111110111100001010010,
    22'b1111111001010001111011,
    22'b1111111010111000010100,
    22'b1111111100001010001111,
    22'b1111111101010001111011,
    22'b1111111101010001111011,
    22'b1111111100111101011100,
    22'b1111111100011110101110,
    22'b1111111011100001010010,
    22'b1111111010111000010100,
    22'b1111111010001111010111,
    22'b1111111001000111101100,
    22'b1111111000000000000000,
    22'b1111110111000010100100,
    22'b1111110110001111010111,
    22'b1111110110000101001000,
    22'b1111110110001111010111,
    22'b1111110110100011110110,
    22'b1111110111010111000011,
    22'b1111110111110101110001,
    22'b1111111000101000111101,
    22'b1111111000101000111101,
    22'b1111111000011110101110,
    22'b1111111000010100011111,
    22'b1111111000000000000000,
    22'b1111110111100001010010,
    22'b1111110111000010100100,
    22'b1111110111001100110011,
    22'b1111110111100001010010,
    22'b1111110111110101110001,
    22'b1111110111110101110001,
    22'b1111110111110101110001,
    22'b1111110111001100110011,
    22'b1111110110011001100110,
    22'b1111110101111010111000,
    22'b1111110101010001111011,
    22'b1111110100111101011100,
    22'b1111110100111101011100,
    22'b1111110100110011001101,
    22'b1111110100101000111101,
    22'b1111110100010100011111,
    22'b1111110100000000000000,
    22'b1111110011100001010010,
    22'b1111110011000010100100,
    22'b1111110010111000010100,
    22'b1111110010111000010100,
    22'b1111110011000010100100,
    22'b1111110011001100110011,
    22'b1111110011100001010010,
    22'b1111110100000000000000,
    22'b1111110100001010001111,
    22'b1111110100111101011100,
    22'b1111110110101110000101,
    22'b1111110110101110000101,
    22'b1111110111001100110011,
    22'b1111110111010111000011,
    22'b1111110111010111000011,
    22'b1111110111001100110011,
    22'b1111110111000010100100,
    22'b1111110111010111000011,
    22'b1111111000011110101110,
    22'b1111110101110000101001,
    22'b1111110001100110011010,
    22'b1111101100011110101110,
    22'b1111100111001100110011,
    22'b1111100010001111010111,
    22'b1111100000111101011100,
    22'b1111100001011100001010,
    22'b1111100011100001010010,
    22'b1111100100101000111101,
    22'b1111100100111101011100,
    22'b1111100100110011001101,
    22'b1111100110100011110110,
    22'b1111101000011110101110,
    22'b1111101011101011100001,
    22'b1111101111110101110001,
    22'b1111110110001111010111,
    22'b1111111001110000101001,
    22'b1111111011110101110001,
    22'b1111111101000111101100,
    22'b1111111101100110011010,
    22'b1111111110011001100110,
    22'b1111111111101011100001,
    22'b0000000010000101001000,
    22'b0000000100000000000000,
    22'b0000000101111010111000,
    22'b0000001100110011001101,
    22'b0000001100011110101110,
    22'b0000001010111000010100,
    22'b0000001000011110101110,
    22'b0000000011100001010010,
    22'b1111111110101110000101,
    22'b1111111001100110011010,
    22'b1111110100101000111101,
    22'b1111101110100011110110,
    22'b1111101010100011110110,
    22'b1111100111101011100001,
    22'b1111100101100110011010,
    22'b1111100100011110101110,
    22'b1111100100110011001101,
    22'b1111100110000101001000,
    22'b1111101000000000000000,
    22'b1111101010111000010100,
    22'b1111101101010001111011,
    22'b1111101111100001010010,
    22'b1111110010011001100110,
    22'b1111110100000000000000,
    22'b1111110101011100001010,
    22'b1111110110011001100110,
    22'b1111110111001100110011,
    22'b1111110111101011100001,
    22'b1111111000001010001111,
    22'b1111111000101000111101,
    22'b1111111001010001111011,
    22'b1111111001110000101001,
    22'b1111111010001111010111,
    22'b1111111010011001100110,
    22'b1111111010001111010111,
    22'b1111111001111010111000,
    22'b1111111001011100001010,
    22'b1111111000111101011100,
    22'b1111111000010100011111,
    22'b1111111000000000000000,
    22'b1111111000000000000000,
    22'b1111111000001010001111,
    22'b1111111000010100011111,
    22'b1111111000010100011111,
    22'b1111111000001010001111,
    22'b1111111000001010001111,
    22'b1111111000101000111101,
    22'b1111111001010001111011,
    22'b1111111001111010111000,
    22'b1111111010100011110110,
    22'b1111111011001100110011,
    22'b1111111011100001010010,
    22'b1111111100000000000000,
    22'b1111111100011110101110,
    22'b1111111101011100001010,
    22'b1111111101111010111000,
    22'b1111111110001111010111,
    22'b1111111110111000010100,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111111100001010010,
    22'b1111111110111000010100,
    22'b1111111110101110000101,
    22'b1111111110101110000101,
    22'b1111111110011001100110,
    22'b1111111101111010111000,
    22'b1111111101100110011010,
    22'b1111111100111101011100,
    22'b1111111011110101110001,
    22'b1111111010011001100110,
    22'b1111111000010100011111,
    22'b1111110110111000010100,
    22'b1111110101110000101001,
    22'b1111110101000111101100,
    22'b1111110101000111101100,
    22'b1111110101010001111011,
    22'b1111110101011100001010,
    22'b1111110101100110011010,
    22'b1111110101100110011010,
    22'b1111110101011100001010,
    22'b1111110101010001111011,
    22'b1111110101010001111011,
    22'b1111110101110000101001,
    22'b1111110101111010111000,
    22'b1111110110000101001000,
    22'b1111110110000101001000,
    22'b1111110110001111010111,
    22'b1111110110000101001000,
    22'b1111110110001111010111,
    22'b1111110110001111010111,
    22'b1111110101111010111000,
    22'b1111110101010001111011,
    22'b1111110100011110101110,
    22'b1111110011110101110001,
    22'b1111110011010111000011,
    22'b1111110010111000010100,
    22'b1111110010011001100110,
    22'b1111110001110000101001,
    22'b1111110000111101011100,
    22'b1111110000011110101110,
    22'b1111110000001010001111,
    22'b1111101111110101110001,
    22'b1111101111100001010010,
    22'b1111101111001100110011,
    22'b1111101111000010100100,
    22'b1111101111001100110011,
    22'b1111101111101011100001,
    22'b1111110000010100011111,
    22'b1111110001000111101100,
    22'b1111110001111010111000,
    22'b1111110011001100110011,
    22'b1111110011110101110001,
    22'b1111110100010100011111,
    22'b1111110100011110101110,
    22'b1111110011100001010010,
    22'b1111110010001111010111,
    22'b1111110001000111101100,
    22'b1111101110001111010111,
    22'b1111101011101011100001,
    22'b1111101001010001111011,
    22'b1111100110100011110110,
    22'b1111100101011100001010,
    22'b1111100101111010111000,
    22'b1111100110100011110110,
    22'b1111101000000000000000,
    22'b1111101001111010111000,
    22'b1111101011001100110011,
    22'b1111101011010111000011,
    22'b1111101011100001010010,
    22'b1111101011101011100001,
    22'b1111101100001010001111,
    22'b1111101100001010001111,
    22'b1111101011101011100001,
    22'b1111101010101110000101,
    22'b1111101001100110011010,
    22'b1111101000101000111101,
    22'b1111100111110101110001,
    22'b1111100111100001010010,
    22'b1111100111000010100100,
    22'b1111100110101110000101,
    22'b1111100110100011110110,
    22'b1111100110011001100110,
    22'b1111100110011001100110,
    22'b1111100110001111010111,
    22'b1111100110000101001000,
    22'b1111100110001111010111,
    22'b1111100110011001100110,
    22'b1111100111010111000011,
    22'b1111101000010100011111,
    22'b1111101001000111101100,
    22'b1111101001111010111000,
    22'b1111101010011001100110,
    22'b1111101011010111000011,
    22'b1111101100010100011111,
    22'b1111101110000101001000,
    22'b1111101110100011110110,
    22'b1111101111010111000011,
    22'b1111110000001010001111,
    22'b1111110001000111101100,
    22'b1111110001111010111000,
    22'b1111110010101110000101,
    22'b1111110011100001010010,
    22'b1111110101000111101100,
    22'b1111110110011001100110,
    22'b1111110111101011100001,
    22'b1111111000110011001101,
    22'b1111111001110000101001,
    22'b1111111010000101001000,
    22'b1111111001111010111000,
    22'b1111111010000101001000,
    22'b1111111010011001100110,
    22'b1111111010111000010100,
    22'b1111111011010111000011,
    22'b1111111011101011100001,
    22'b1111111011110101110001,
    22'b1111111011110101110001,
    22'b1111111011110101110001,
    22'b1111111011100001010010,
    22'b1111111011001100110011,
    22'b1111111010111000010100,
    22'b1111111010101110000101,
    22'b1111111010011001100110,
    22'b1111111010000101001000,
    22'b1111111001110000101001,
    22'b1111111000111101011100,
    22'b1111110111001100110011,
    22'b1111110110001111010111,
    22'b1111110101100110011010,
    22'b1111110100001010001111,
    22'b1111110011000010100100,
    22'b1111110010101110000101,
    22'b1111110100001010001111,
    22'b1111110011001100110011,
    22'b1111110101011100001010,
    22'b1111110111000010100100,
    22'b1111111000010100011111,
    22'b1111111010001111010111,
    22'b1111111011100001010010,
    22'b1111111100101000111101,
    22'b1111111101011100001010,
    22'b1111111111001100110011,
    22'b0000000000010100011111,
    22'b0000000001010001111011,
    22'b0000000010111000010100,
    22'b0000000100011110101110,
    22'b0000000101111010111000,
    22'b0000000110111000010100,
    22'b0000001000001010001111,
    22'b0000001001011100001010,
    22'b0000001011000010100100,
    22'b0000001100111101011100,
    22'b0000001111110101110001,
    22'b0000010001111010111000,
    22'b0000010011101011100001,
    22'b0000010101010001111011,
    22'b0000010111001100110011,
    22'b0000011000010100011111,
    22'b0000011001000111101100,
    22'b0000011100010100011111,
    22'b0000011101110000101001,
    22'b0000011111101011100001,
    22'b0000100001111010111000,
    22'b0000100100110011001101,
    22'b0000100111000010100100,
    22'b0000101001000111101100,
    22'b0000101011010111000011,
    22'b0000101100101000111101,
    22'b0000101101100110011010,
    22'b0000101110001111010111,
    22'b0000101110100011110110,
    22'b0000101110100011110110,
    22'b0000101110001111010111,
    22'b0000101110000101001000,
    22'b0000101101111010111000,
    22'b0000101101011100001010,
    22'b0000101101010001111011,
    22'b0000101101011100001010,
    22'b0000101110100011110110,
    22'b0000101111110101110001,
    22'b0000110000110011001101,
    22'b0000110000111101011100,
    22'b0000110000010100011111,
    22'b0000101111001100110011,
    22'b0000101110000101001000,
    22'b0000101101100110011010,
    22'b0000101101011100001010,
    22'b0000101101011100001010,
    22'b0000101101100110011010,
    22'b0000101101110000101001,
    22'b0000101101111010111000,
    22'b0000101110000101001000,
    22'b0000101110000101001000,
    22'b0000101101011100001010,
    22'b0000101100101000111101,
    22'b0000101011101011100001,
    22'b0000101010011001100110,
    22'b0000101000010100011111,
    22'b0000100110101110000101,
    22'b0000100101000111101100,
    22'b0000100011010111000011,
    22'b0000100001011100001010,
    22'b0000100000000000000000,
    22'b0000011110011001100110,
    22'b0000011100101000111101,
    22'b0000011001110000101001,
    22'b0000010111101011100001,
    22'b0000010101100110011010,
    22'b0000010011110101110001,
    22'b0000010001110000101001,
    22'b0000010000010100011111,
    22'b0000001110111000010100,
    22'b0000001101100110011010,
    22'b0000001100010100011111,
    22'b0000001010011001100110,
    22'b0000001000111101011100,
    22'b0000000111101011100001,
    22'b0000000110100011110110,
    22'b0000000101010001111011,
    22'b0000000100110011001101,
    22'b0000000100010100011111,
    22'b0000000100001010001111,
    22'b0000000100000000000000,
    22'b0000000011101011100001,
    22'b0000000011010111000011,
    22'b0000000011000010100100,
    22'b0000000011000010100100,
    22'b0000000011010111000011,
    22'b0000000011101011100001,
    22'b0000000100001010001111,
    22'b0000000100110011001101,
    22'b0000000101011100001010,
    22'b0000001100000000000000,
    22'b0000001011100001010010,
    22'b0000001000101000111101,
    22'b0000000000110011001101,
    22'b1111111010011001100110,
    22'b1111110011110101110001,
    22'b1111101110101110000101,
    22'b1111101001111010111000,
    22'b1111100111000010100100,
    22'b1111100101011100001010,
    22'b1111100100111101011100,
    22'b1111100100110011001101,
    22'b1111100101000111101100,
    22'b1111100101011100001010,
    22'b1111100101110000101001,
    22'b1111100110001111010111,
    22'b1111100111001100110011,
    22'b1111101000001010001111,
    22'b1111101001000111101100,
    22'b1111101010011001100110,
    22'b1111101100010100011111,
    22'b1111101101111010111000,
    22'b1111101111101011100001,
    22'b1111110001011100001010,
    22'b1111110011110101110001,
    22'b1111110101100110011010,
    22'b1111110111001100110011,
    22'b1111111000110011001101,
    22'b1111111010111000010100,
    22'b1111111100001010001111,
    22'b1111111101000111101100,
    22'b1111111101110000101001,
    22'b1111111101111010111000,
    22'b1111111101111010111000,
    22'b1111111101110000101001,
    22'b1111111101110000101001,
    22'b1111111110000101001000,
    22'b1111111110011001100110,
    22'b1111111110111000010100,
    22'b1111111111010111000011,
    22'b1111111111101011100001,
    22'b1111111111101011100001,
    22'b1111111111010111000011,
    22'b1111111110011001100110,
    22'b1111111100011110101110,
    22'b1111111011000010100100,
    22'b1111111001011100001010,
    22'b1111111000001010001111,
    22'b1111110110111000010100,
    22'b1111110110000101001000,
    22'b1111110101110000101001,
    22'b1111110101011100001010,
    22'b1111110101010001111011,
    22'b1111110101000111101100,
    22'b1111110100111101011100,
    22'b1111110100010100011111,
    22'b1111110011010111000011,
    22'b1111110010100011110110,
    22'b1111110001100110011010,
    22'b1111101111010111000011,
    22'b1111101111010111000011,
    22'b1111110000000000000000,
    22'b1111110000111101011100,
    22'b1111110010100011110110,
    22'b1111110011110101110001,
    22'b1111110101000111101100,
    22'b1111110110001111010111,
    22'b1111110111110101110001,
    22'b1111111001000111101100,
    22'b1111111010000101001000,
    22'b1111111010111000010100,
    22'b1111111011100001010010,
    22'b1111111100001010001111,
    22'b1111111100010100011111,
    22'b1111111100001010001111,
    22'b1111111100000000000000,
    22'b1111111011100001010010,
    22'b1111111010101110000101,
    22'b1111111010000101001000,
    22'b1111111001000111101100,
    22'b1111111000000000000000,
    22'b1111110111000010100100,
    22'b1111110110001111010111,
    22'b1111110101000111101100,
    22'b1111110100011110101110,
    22'b1111110011101011100001,
    22'b1111110011000010100100,
    22'b1111110010100011110110,
    22'b1111110010011001100110,
    22'b1111110010011001100110,
    22'b1111110010101110000101,
    22'b1111110011100001010010,
    22'b1111110100001010001111,
    22'b1111110100110011001101,
    22'b1111110101100110011010,
    22'b1111110110100011110110,
    22'b1111110111010111000011,
    22'b1111111000001010001111,
    22'b1111111001000111101100,
    22'b1111111010001111010111,
    22'b1111111011000010100100,
    22'b1111111100000000000000,
    22'b1111111100110011001101,
    22'b1111111101111010111000,
    22'b1111111110101110000101,
    22'b1111111111010111000011,
    22'b1111111111110101110001,
    22'b0000000001010001111011,
    22'b0000000001011100001010,
    22'b0000000001100110011010,
    22'b0000000001000111101100,
    22'b0000000000011110101110,
    22'b0000000001000111101100,
    22'b0000000010000101001000,
    22'b0000000011100001010010,
    22'b0000000101011100001010,
    22'b0000000101100110011010,
    22'b0000000111100001010010,
    22'b0000010001011100001010,
    22'b0000010100001010001111,
    22'b0000010000000000000000,
    22'b0000001100011110101110,
    22'b0000000100011110101110,
    22'b1111111111100001010010,
    22'b1111111101110000101001,
    22'b1111111100011110101110,
    22'b1111111001010001111011,
    22'b1111111000000000000000,
    22'b1111111000001010001111,
    22'b1111111010011001100110,
    22'b1111111101011100001010,
    22'b0000000000110011001101,
    22'b0000000011001100110011,
    22'b0000000100110011001101,
    22'b0000000100111101011100,
    22'b0000000100110011001101,
    22'b0000000100110011001101,
    22'b0000000100111101011100,
    22'b0000000100110011001101,
    22'b0000000100011110101110,
    22'b0000000011101011100001,
    22'b0000000010011001100110,
    22'b0000000001010001111011,
    22'b0000000000010100011111,
    22'b1111111111110101110001,
    22'b0000000000000000000000,
    22'b0000000000000000000000,
    22'b0000000000001010001111,
    22'b0000000000010100011111,
    22'b0000000000011110101110,
    22'b0000000000110011001101,
    22'b0000000001010001111011,
    22'b0000000001111010111000,
    22'b0000000010001111010111,
    22'b0000000010100011110110,
    22'b0000000010011001100110,
    22'b0000000001110000101001,
    22'b0000000001000111101100,
    22'b0000000000010100011111,
    22'b1111111111100001010010,
    22'b1111111110101110000101,
    22'b1111111110000101001000,
    22'b1111111101100110011010,
    22'b1111111101011100001010,
    22'b1111111101010001111011,
    22'b1111111101010001111011,
    22'b1111111101010001111011,
    22'b1111111101011100001010,
    22'b1111111101110000101001,
    22'b1111111101111010111000,
    22'b1111111101111010111000,
    22'b1111111101100110011010,
    22'b1111111101000111101100,
    22'b1111111100011110101110,
    22'b1111111011110101110001,
    22'b1111111011001100110011,
    22'b1111111010101110000101,
    22'b1111111010001111010111,
    22'b1111111001111010111000,
    22'b1111111001110000101001,
    22'b1111111001110000101001,
    22'b1111111001111010111000,
    22'b1111111010000101001000,
    22'b1111111010011001100110,
    22'b1111111010111000010100,
    22'b1111111010011001100110,
    22'b1111111001010001111011,
    22'b1111111000000000000000,
    22'b1111110111000010100100,
    22'b1111110110000101001000,
    22'b1111110101010001111011,
    22'b1111110101010001111011,
    22'b1111110101100110011010,
    22'b1111110110001111010111,
    22'b1111110111000010100100,
    22'b1111110111110101110001,
    22'b1111111001000111101100,
    22'b1111111011000010100100,
    22'b1111111100110011001101,
    22'b1111111110101110000101,
    22'b0000000000011110101110,
    22'b0000000010000101001000,
    22'b0000000011100001010010,
    22'b0000000100011110101110,
    22'b0000000101010001111011,
    22'b0000000110000101001000,
    22'b0000000110101110000101,
    22'b0000000111001100110011,
    22'b0000000111010111000011,
    22'b0000000111100001010010,
    22'b0000000111101011100001,
    22'b0000001000000000000000,
    22'b0000001000010100011111,
    22'b0000001000011110101110,
    22'b0000001000010100011111,
    22'b0000001000000000000000,
    22'b0000000111010111000011,
    22'b0000000110101110000101,
    22'b0000000110000101001000,
    22'b0000000101011100001010,
    22'b0000000100110011001101,
    22'b0000000100000000000000,
    22'b0000000011110101110001,
    22'b0000000100000000000000,
    22'b0000000100110011001101,
    22'b0000000110001111010111,
    22'b0000000111100001010010,
    22'b0000001000111101011100,
    22'b0000001010000101001000,
    22'b0000001011001100110011,
    22'b0000001100000000000000,
    22'b0000001100101000111101,
    22'b0000001100111101011100,
    22'b0000001101000111101100,
    22'b0000001101000111101100,
    22'b0000001100101000111101,
    22'b0000001011110101110001,
    22'b0000001011000010100100,
    22'b0000001010000101001000,
    22'b0000001000110011001101,
    22'b0000001000000000000000,
    22'b0000000110101110000101,
    22'b0000000101111010111000,
    22'b0000000100011110101110,
    22'b0000000011101011100001,
    22'b0000000010100011110110,
    22'b0000000001111010111000,
    22'b0000000001010001111011,
    22'b0000000000110011001101,
    22'b0000000001000111101100,
    22'b0000000001111010111000,
    22'b0000000011000010100100,
    22'b0000000100110011001101,
    22'b0000000110001111010111,
    22'b0000000111100001010010,
    22'b0000001000101000111101,
    22'b0000001001100110011010,
    22'b0000001011000010100100,
    22'b0000001011101011100001,
    22'b0000001100010100011111,
    22'b0000001100110011001101,
    22'b0000001101010001111011,
    22'b0000001110100011110110,
    22'b0000001110111000010100,
    22'b0000001110101110000101,
    22'b0000001110101110000101,
    22'b0000001110101110000101,
    22'b0000001110001111010111,
    22'b0000001101111010111000,
    22'b0000001101010001111011,
    22'b0000001100010100011111,
    22'b0000001011000010100100,
    22'b0000001010001111010111,
    22'b0000001001110000101001,
    22'b0000001001110000101001,
    22'b0000001010100011110110,
    22'b0000001011010111000011,
    22'b0000001011110101110001,
    22'b0000001011101011100001,
    22'b0000001011000010100100,
    22'b0000001010011001100110,
    22'b0000001010000101001000,
    22'b0000001010011001100110,
    22'b0000001011010111000011,
    22'b0000001101010001111011,
    22'b0000001110000101001000,
    22'b0000001110000101001000,
    22'b0000001101110000101001,
    22'b0000001101000111101100,
    22'b0000001100110011001101,
    22'b0000001011101011100001,
    22'b0000001010000101001000,
    22'b0000001000011110101110,
    22'b0000000110011001100110,
    22'b0000000101000111101100,
    22'b0000000011110101110001,
    22'b0000000011000010100100,
    22'b0000000010100011110110,
    22'b0000000010001111010111,
    22'b0000000010011001100110,
    22'b0000000010011001100110,
    22'b0000000010101110000101,
    22'b0000000011001100110011,
    22'b0000000011010111000011,
    22'b0000000011100001010010,
    22'b0000000011101011100001,
    22'b0000000011100001010010,
    22'b0000000011001100110011,
    22'b0000000011000010100100,
    22'b0000000010111000010100,
    22'b0000000010100011110110,
    22'b0000000001100110011010,
    22'b0000000000101000111101,
    22'b1111111111101011100001,
    22'b1111111110101110000101,
    22'b1111111110000101001000,
    22'b1111111101110000101001,
    22'b1111111101111010111000,
    22'b1111111110001111010111,
    22'b1111111110011001100110,
    22'b1111111110000101001000,
    22'b1111111101110000101001,
    22'b1111111101100110011010,
    22'b1111111101111010111000,
    22'b1111111110011001100110,
    22'b1111111111010111000011,
    22'b0000000000001010001111,
    22'b0000000000110011001101,
    22'b0000000001000111101100,
    22'b0000000001100110011010,
    22'b0000000001111010111000,
    22'b0000000001111010111000,
    22'b1111111011101011100001,
    22'b1111110010011001100110,
    22'b1111011100001010001111,
    22'b1111011110101110000101,
    22'b1111100001000111101100,
    22'b1111100011010111000011,
    22'b1111100100010100011111,
    22'b1111100100111101011100,
    22'b1111100101010001111011,
    22'b1111100101100110011010,
    22'b1111100110000101001000,
    22'b1111100110100011110110,
    22'b1111100111010111000011,
    22'b1111101000010100011111,
    22'b1111101001110000101001,
    22'b1111101010101110000101,
    22'b1111101011100001010010,
    22'b1111101011110101110001,
    22'b1111101011110101110001,
    22'b1111101011010111000011,
    22'b1111101010101110000101,
    22'b1111101001110000101001,
    22'b1111101000101000111101,
    22'b1111100111110101110001,
    22'b1111100111001100110011,
    22'b1111100110111000010100,
    22'b1111100111000010100100,
    22'b1111100111101011100001,
    22'b1111101000110011001101,
    22'b1111101010011001100110,
    22'b1111101100001010001111,
    22'b1111101110001111010111,
    22'b1111101111001100110011,
    22'b1111110000010100011111,
    22'b1111110001000111101100,
    22'b1111110010000101001000,
    22'b1111110011000010100100,
    22'b1111110100001010001111,
    22'b1111110101011100001010,
    22'b1111110111101011100001,
    22'b1111111001100110011010,
    22'b1111111011010111000011,
    22'b1111111100111101011100,
    22'b1111111110111000010100,
    22'b0000000000000000000000,
    22'b0000000001000111101100,
    22'b0000000010001111010111,
    22'b0000000011101011100001,
    22'b0000000100110011001101,
    22'b0000000101100110011010,
    22'b0000000110001111010111,
    22'b0000000110100011110110,
    22'b0000000110100011110110,
    22'b0000000110001111010111,
    22'b0000000101111010111000,
    22'b0000000101011100001010,
    22'b0000000100110011001101,
    22'b0000000100001010001111,
    22'b0000000011100001010010,
    22'b0000000010111000010100,
    22'b0000000001100110011010,
    22'b0000000000011110101110,
    22'b1111111111100001010010,
    22'b1111111110100011110110,
    22'b1111111101011100001010,
    22'b1111111100000000000000,
    22'b1111111011000010100100,
    22'b1111111010000101001000,
    22'b1111111001010001111011,
    22'b1111111000010100011111,
    22'b1111110111110101110001,
    22'b1111110111100001010010,
    22'b1111110111000010100100,
    22'b1111110110001111010111,
    22'b1111110101100110011010,
    22'b1111110100111101011100,
    22'b1111110100111101011100,
    22'b1111110101100110011010,
    22'b1111110110100011110110,
    22'b1111110111101011100001,
    22'b1111111011100001010010,
    22'b1111111100000000000000,
    22'b1111111100000000000000,
    22'b1111111011101011100001,
    22'b1111111010011001100110,
    22'b1111111000111101011100,
    22'b1111110111100001010010,
    22'b1111110101111010111000,
    22'b1111110100000000000000,
    22'b1111110010011001100110,
    22'b1111110000101000111101,
    22'b1111101110111000010100,
    22'b1111101100110011001101,
    22'b1111101011101011100001,
    22'b1111101010111000010100,
    22'b1111101010100011110110,
    22'b1111101010100011110110,
    22'b1111101010101110000101,
    22'b1111101011000010100100,
    22'b1111101011001100110011,
    22'b1111101011010111000011,
    22'b1111101011100001010010,
    22'b1111101011100001010010,
    22'b1111101011110101110001,
    22'b1111101100001010001111,
    22'b1111101100101000111101,
    22'b1111101101010001111011,
    22'b1111101110011001100110,
    22'b1111101111001100110011,
    22'b1111101111110101110001,
    22'b1111110000011110101110,
    22'b1111110001010001111011,
    22'b1111110001100110011010,
    22'b1111110001110000101001,
    22'b1111110001100110011010,
    22'b1111110000111101011100,
    22'b1111110000001010001111,
    22'b1111101111010111000011,
    22'b1111101111100001010010,
    22'b1111110000001010001111,
    22'b1111110000010100011111,
    22'b1111110000000000000000,
    22'b1111101110111000010100,
    22'b1111101110001111010111,
    22'b1111101101110000101001,
    22'b1111101101110000101001,
    22'b1111101110100011110110,
    22'b1111101111100001010010,
    22'b1111110000110011001101,
    22'b1111110010001111010111,
    22'b1111110100000000000000,
    22'b1111110101000111101100,
    22'b1111110101111010111000,
    22'b1111110110000101001000,
    22'b1111110101100110011010,
    22'b1111110100111101011100,
    22'b1111110100000000000000,
    22'b1111110011001100110011,
    22'b1111110010101110000101,
    22'b1111110010011001100110,
    22'b1111110010000101001000,
    22'b1111110001110000101001,
    22'b1111110001100110011010,
    22'b1111110001100110011010,
    22'b1111110010000101001000,
    22'b1111110010100011110110,
    22'b1111110011000010100100,
    22'b1111110011100001010010,
    22'b1111110011110101110001,
    22'b1111110011110101110001,
    22'b1111110011101011100001,
    22'b1111110011010111000011,
    22'b1111110010111000010100,
    22'b1111110010101110000101,
    22'b1111110010100011110110,
    22'b1111110000000000000000,
    22'b1111101111100001010010,
    22'b1111101111010111000011,
    22'b1111101110111000010100,
    22'b1111101110101110000101,
    22'b1111101110101110000101,
    22'b1111101111000010100100,
    22'b1111110000000000000000,
    22'b1111110001000111101100,
    22'b1111110010000101001000,
    22'b1111110010101110000101,
    22'b1111110010111000010100,
    22'b1111110010001111010111,
    22'b1111110001010001111011,
    22'b1111101111110101110001,
    22'b1111101110100011110110,
    22'b1111101101011100001010,
    22'b1111101100010100011111,
    22'b1111101011000010100100,
    22'b1111101010001111010111,
    22'b1111101001100110011010,
    22'b1111101001000111101100,
    22'b1111101000111101011100,
    22'b1111101000101000111101,
    22'b1111101000110011001101,
    22'b1111101000111101011100,
    22'b1111101001000111101100,
    22'b1111101001010001111011,
    22'b1111101001000111101100,
    22'b1111101001000111101100,
    22'b1111101001000111101100,
    22'b1111101000111101011100,
    22'b1111101001010001111011,
    22'b1111101001110000101001,
    22'b1111101010000101001000,
    22'b1111101010100011110110,
    22'b1111101010111000010100,
    22'b1111101011001100110011,
    22'b1111101011101011100001,
    22'b1111101100010100011111,
    22'b1111101100101000111101,
    22'b1111101100111101011100,
    22'b1111101101010001111011,
    22'b1111101101110000101001,
    22'b1111101110011001100110,
    22'b1111101111001100110011,
    22'b1111110000010100011111,
    22'b1111110001010001111011,
    22'b1111110010000101001000,
    22'b1111110010111000010100,
    22'b1111110100000000000000,
    22'b1111110100101000111101,
    22'b1111110101000111101100,
    22'b1111110101011100001010,
    22'b1111110101011100001010,
    22'b1111110101010001111011,
    22'b1111110100111101011100,
    22'b1111110100011110101110,
    22'b1111110100001010001111,
    22'b1111110011101011100001,
    22'b1111110010111000010100,
    22'b1111110001100110011010,
    22'b1111101111010111000011,
    22'b1111101111100001010010,
    22'b1111101111001100110011,
    22'b1111101110100011110110,
    22'b1111101110000101001000,
    22'b1111101101011100001010,
    22'b1111101101000111101100,
    22'b1111101100111101011100,
    22'b1111101100111101011100,
    22'b1111101100101000111101,
    22'b1111101100001010001111,
    22'b1111101011100001010010,
    22'b1111101010111000010100,
    22'b1111101010001111010111,
    22'b1111101010000101001000,
    22'b1111101010000101001000,
    22'b1111101010001111010111,
    22'b1111101010011001100110,
    22'b1111101010100011110110,
    22'b1111101010100011110110,
    22'b1111101010101110000101,
    22'b1111101010101110000101,
    22'b1111101010101110000101,
    22'b1111101010101110000101,
    22'b1111101010100011110110,
    22'b1111101010011001100110,
    22'b1111101010001111010111,
    22'b1111101010000101001000,
    22'b1111101010001111010111,
    22'b1111101010100011110110,
    22'b1111101011000010100100,
    22'b1111101001011100001010,
    22'b1111100111110101110001,
    22'b1111100101110000101001,
    22'b1111100010101110000101,
    22'b1111100000000000000000,
    22'b1111011101100110011010,
    22'b1111011010011001100110,
    22'b1111011000011110101110,
    22'b1111010111000010100100,
    22'b1111010101110000101001,
    22'b1111010100011110101110,
    22'b1111010011101011100001,
    22'b1111010011000010100100,
    22'b1111010010111000010100,
    22'b1111010011001100110011,
    22'b1111010100001010001111,
    22'b1111010101110000101001,
    22'b1111011000010100011111,
    22'b1111011010101110000101,
    22'b1111011101000111101100,
    22'b1111011111101011100001,
    22'b1111100010111000010100,
    22'b1111100100101000111101,
    22'b1111100101111010111000,
    22'b1111100110100011110110,
    22'b1111100110100011110110,
    22'b1111100110000101001000,
    22'b1111100101011100001010,
    22'b1111100101000111101100,
    22'b1111100101000111101100,
    22'b1111101001010001111011,
    22'b1111101010011001100110,
    22'b1111101010011001100110,
    22'b1111101001011100001010,
    22'b1111100110101110000101,
    22'b1111100100000000000000,
    22'b1111100000110011001101,
    22'b1111011101011100001010,
    22'b1111011001000111101100,
    22'b1111010101111010111000,
    22'b1111010010101110000101,
    22'b1111001111101011100001,
    22'b1111001100110011001101,
    22'b1111001011010111000011,
    22'b1111001011000010100100,
    22'b1111001100000000000000,
    22'b1111001101010001111011,
    22'b1111001111000010100100,
    22'b1111010000111101011100,
    22'b1111010011100001010010,
    22'b1111010101110000101001,
    22'b1111010111110101110001,
    22'b1111011010000101001000,
    22'b1111011011010111000011,
    22'b1111011100001010001111,
    22'b1111011100101000111101,
    22'b1111011100111101011100,
    22'b1111011101100110011010,
    22'b1111011110001111010111,
    22'b1111011111000010100100,
    22'b1111100000101000111101,
    22'b1111100010100011110110,
    22'b1111101111000010100100,
    22'b1111110010100011110110,
    22'b1111110100010100011111,
    22'b1111110101010001111011,
    22'b1111110101100110011010,
    22'b1111110101010001111011,
    22'b1111110100101000111101,
    22'b1111110100000000000000,
    22'b1111110011001100110011,
    22'b1111110010100011110110,
    22'b1111110001111010111000,
    22'b1111110001000111101100,
    22'b1111110000000000000000,
    22'b1111101111010111000011,
    22'b1111101111000010100100,
    22'b1111101111000010100100,
    22'b1111101111100001010010,
    22'b1111110000001010001111,
    22'b1111110000110011001101,
    22'b1111110001011100001010,
    22'b1111110001111010111000,
    22'b1111110010001111010111,
    22'b1111110010011001100110,
    22'b1111110010100011110110,
    22'b1111110010001111010111,
    22'b1111110001011100001010,
    22'b1111101110111000010100,
    22'b1111101101000111101100,
    22'b1111100101111010111000,
    22'b1111100100111101011100,
    22'b1111100100011110101110,
    22'b1111100100010100011111,
    22'b1111100100000000000000,
    22'b1111100100000000000000,
    22'b1111100100001010001111,
    22'b1111100100001010001111,
    22'b1111100100011110101110,
    22'b1111100100010100011111,
    22'b1111100011101011100001,
    22'b1111100010101110000101,
    22'b1111100000000000000000,
    22'b1111011101010001111011,
    22'b1111011010011001100110,
    22'b1111010110111000010100,
    22'b1111010101000111101100,
    22'b1111010100000000000000,
    22'b1111010010101110000101,
    22'b1111010010100011110110,
    22'b1111010010000101001000,
    22'b1111010010101110000101,
    22'b1111010011101011100001,
    22'b1111010101010001111011,
    22'b1111010111010111000011,
    22'b1111011000101000111101,
    22'b1111011001100110011010,
    22'b1111011010011001100110,
    22'b1111011010000101001000,
    22'b1111011010001111010111,
    22'b1111011100111101011100,
    22'b1111011101000111101100,
    22'b1111011101010001111011,
    22'b1111011101010001111011,
    22'b1111011100101000111101,
    22'b1111011100101000111101,
    22'b1111011100101000111101,
    22'b1111011100011110101110,
    22'b1111011100011110101110,
    22'b1111011101010001111011,
    22'b1111011110001111010111,
    22'b1111011111100001010010,
    22'b1111100000101000111101,
    22'b1111100001110000101001,
    22'b1111100010101110000101,
    22'b1111100100010100011111,
    22'b1111100101011100001010,
    22'b1111100110111000010100,
    22'b1111101000000000000000,
    22'b1111101001010001111011,
    22'b1111101010100011110110,
    22'b1111101011101011100001,
    22'b1111101100101000111101,
    22'b1111101100111101011100,
    22'b1111101100001010001111,
    22'b1111101011110101110001,
    22'b1111101100000000000000,
    22'b1111101100011110101110,
    22'b1111101101000111101100,
    22'b1111101110101110000101,
    22'b1111110001111010111000,
    22'b1111101111101011100001,
    22'b1111101110011001100110,
    22'b1111101110011001100110,
    22'b1111110000011110101110,
    22'b1111110010100011110110,
    22'b1111110100101000111101,
    22'b1111110110100011110110,
    22'b1111110111110101110001,
    22'b1111111000001010001111,
    22'b1111111001011100001010,
    22'b1111111010001111010111,
    22'b1111111010001111010111,
    22'b1111111001110000101001,
    22'b1111111000101000111101,
    22'b1111110111100001010010,
    22'b1111110110001111010111,
    22'b1111110101110000101001,
    22'b1111110110000101001000,
    22'b1111110110111000010100,
    22'b1111110111100001010010,
    22'b1111110111010111000011,
    22'b1111110111001100110011,
    22'b1111110110111000010100,
    22'b1111110110111000010100,
    22'b1111110110101110000101,
    22'b1111110110111000010100,
    22'b1111110110111000010100,
    22'b1111110110111000010100,
    22'b1111110111101011100001,
    22'b1111111000110011001101,
    22'b1111111101011100001010,
    22'b1111111101111010111000,
    22'b1111111110100011110110,
    22'b1111111111100001010010,
    22'b0000000000000000000000,
    22'b0000000000011110101110,
    22'b0000000000111101011100,
    22'b0000000000111101011100,
    22'b0000000000011110101110,
    22'b1111111111110101110001,
    22'b1111111111010111000011,
    22'b1111111110101110000101,
    22'b1111111110011001100110,
    22'b1111111110100011110110,
    22'b1111111110101110000101,
    22'b1111111110111000010100,
    22'b1111111111001100110011,
    22'b1111111111101011100001,
    22'b0000000000010100011111,
    22'b0000000000110011001101,
    22'b0000000000011110101110,
    22'b1111111111110101110001,
    22'b1111111111000010100100,
    22'b1111111101100110011010,
    22'b1111111100110011001101,
    22'b1111111100001010001111,
    22'b1111111100000000000000,
    22'b1111111011110101110001,
    22'b1111111011100001010010,
    22'b1111111011010111000011,
    22'b1111111011001100110011,
    22'b1111111010111000010100,
    22'b1111111010101110000101,
    22'b1111111010100011110110,
    22'b1111111010100011110110,
    22'b1111111010100011110110,
    22'b1111111010100011110110,
    22'b1111111011000010100100,
    22'b1111111011110101110001,
    22'b1111111101100110011010,
    22'b1111111111010111000011,
    22'b0000000000101000111101,
    22'b0000000001011100001010,
    22'b0000000001111010111000,
    22'b0000000001100110011010,
    22'b0000000001110000101001,
    22'b0000000001011100001010,
    22'b0000000001011100001010,
    22'b0000000001000111101100,
    22'b0000000000011110101110,
    22'b1111111111101011100001,
    22'b1111111110101110000101,
    22'b1111111110001111010111,
    22'b1111111110001111010111,
    22'b1111111110001111010111,
    22'b1111111110101110000101,
    22'b1111111111001100110011,
    22'b1111111111100001010010,
    22'b0000000000000000000000,
    22'b0000000000011110101110,
    22'b0000000001000111101100,
    22'b0000000001011100001010,
    22'b0000000010000101001000,
    22'b0000000011001100110011,
    22'b0000000011110101110001,
    22'b0000000100101000111101,
    22'b0000000101100110011010,
    22'b0000000111000010100100,
    22'b0000001000001010001111,
    22'b0000001001011100001010,
    22'b0000001010101110000101,
    22'b0000001100101000111101,
    22'b0000001110011001100110,
    22'b0000010101111010111000,
    22'b0000010110011001100110,
    22'b0000010101110000101001,
    22'b0000010011101011100001,
    22'b0000010000101000111101,
    22'b0000001100110011001101,
    22'b0000000111101011100001,
    22'b0000000100010100011111,
    22'b0000000001111010111000,
    22'b0000000000011110101110,
    22'b0000000000000000000000,
    22'b0000000000101000111101,
    22'b0000000001110000101001,
    22'b0000000011001100110011,
    22'b0000000100110011001101,
    22'b0000000101111010111000,
    22'b0000000111001100110011,
    22'b0000001000101000111101,
    22'b0000001010100011110110,
    22'b0000001100001010001111,
    22'b0000001101011100001010,
    22'b0000001110100011110110,
    22'b0000001111101011100001,
    22'b0000010000011110101110,
    22'b0000010000111101011100,
    22'b0000010001011100001010,
    22'b0000010001111010111000,
    22'b0000010010011001100110,
    22'b0000010010100011110110,
    22'b0000010010101110000101,
    22'b0000010010101110000101,
    22'b0000010010100011110110,
    22'b0000010010100011110110,
    22'b0000010010100011110110,
    22'b0000010010101110000101,
    22'b0000010010111000010100,
    22'b0000010011000010100100,
    22'b0000010011001100110011,
    22'b0000010011000010100100,
    22'b0000010000000000000000,
    22'b0000001111000010100100,
    22'b0000001110000101001000,
    22'b0000001100111101011100,
    22'b0000001100010100011111,
    22'b0000001011101011100001,
    22'b0000001011001100110011,
    22'b0000001010111000010100,
    22'b0000001010101110000101,
    22'b0000001010111000010100,
    22'b0000001011000010100100,
    22'b0000001011010111000011,
    22'b0000001011110101110001,
    22'b0000001100010100011111,
    22'b0000001100111101011100,
    22'b0000001101100110011010,
    22'b0000001110011001100110,
    22'b0000001111100001010010,
    22'b0000010001011100001010,
    22'b0000010011010111000011,
    22'b0000010101010001111011,
    22'b0000010111001100110011,
    22'b0000011001111010111000,
    22'b0000011011101011100001,
    22'b0000011101011100001010,
    22'b0000011111000010100100,
    22'b0000100001010001111011,
    22'b0000100010111000010100,
    22'b0000100100011110101110,
    22'b0000100110001111010111,
    22'b0000101000011110101110,
    22'b0000101010000101001000,
    22'b0000101011101011100001,
    22'b0000101101100110011010,
    22'b0000110000001010001111,
    22'b0000110010001111010111,
    22'b0000110100001010001111,
    22'b0000110110011001100110,
    22'b0000110111101011100001,
    22'b0000111000101000111101,
    22'b0000111001011100001010,
    22'b0000111001111010111000,
    22'b0000111001011100001010,
    22'b0000111000101000111101,
    22'b0000110111100001010010,
    22'b0000110110101110000101,
    22'b0000110101110000101001,
    22'b0000110100101000111101,
    22'b0000110010111000010100,
    22'b0000110001110000101001,
    22'b0000110000101000111101,
    22'b0000101111110101110001,
    22'b0000101111000010100100,
    22'b0000101110111000010100,
    22'b0000101110101110000101,
    22'b0000101111000010100100,
    22'b0000110000000000000000,
    22'b0000110001000111101100,
    22'b0000110010011001100110,
    22'b0000110100001010001111,
    22'b0000110110100011110110,
    22'b0000111000010100011111,
    22'b0000111001110000101001,
    22'b0000111010101110000101,
    22'b0000111011100001010010,
    22'b0000111011101011100001,
    22'b0000111011100001010010,
    22'b0000111011001100110011,
    22'b0000111010101110000101,
    22'b0000111010011001100110,
    22'b0000111010000101001000,
    22'b0000111001110000101001,
    22'b0000111001100110011010,
    22'b0000111001111010111000,
    22'b0000111010001111010111,
    22'b0000111010100011110110,
    22'b0000111010111000010100,
    22'b0000111010111000010100,
    22'b0000111010111000010100,
    22'b0000111010100011110110,
    22'b0000111001111010111000,
    22'b0000111001000111101100,
    22'b0000111000000000000000,
    22'b0000110110101110000101,
    22'b0000110100111101011100,
    22'b0000110010011001100110,
    22'b0000110000011110101110,
    22'b0000101110100011110110,
    22'b0000101100111101011100,
    22'b0000101011001100110011,
    22'b0000101010011001100110,
    22'b0000101001111010111000,
    22'b0000101001100110011010,
    22'b0000101001000111101100,
    22'b0000101001011100001010,
    22'b0000101010101110000101,
    22'b0000101100011110101110,
    22'b0000101110011001100110,
    22'b0000110010101110000101,
    22'b0000110011101011100001,
    22'b0000110100110011001101,
    22'b0000110101011100001010,
    22'b0000110101111010111000,
    22'b0000110110001111010111,
    22'b0000110101111010111000,
    22'b0000110101010001111011,
    22'b0000110100001010001111,
    22'b0000110010101110000101,
    22'b0000110000111101011100,
    22'b0000101110001111010111,
    22'b0000101100000000000000,
    22'b0000101001100110011010,
    22'b0000100111001100110011,
    22'b0000100100010100011111,
    22'b0000100010100011110110,
    22'b0000100001010001111011,
    22'b0000100000010100011111,
    22'b0000011111100001010010,
    22'b0000011110101110000101,
    22'b0000011110000101001000,
    22'b0000011101010001111011,
    22'b0000011100010100011111,
    22'b0000011011010111000011,
    22'b0000011010000101001000,
    22'b0000011000010100011111,
    22'b0000010110000101001000,
    22'b0000010010111000010100,
    22'b0000010001000111101100,
    22'b0000010000001010001111,
    22'b0000010000000000000000,
    22'b0000010000011110101110,
    22'b0000010010000101001000,
    22'b0000010011101011100001,
    22'b0000010101010001111011,
    22'b0000010111000010100100,
    22'b0000011001000111101100,
    22'b0000011010100011110110,
    22'b0000011100000000000000,
    22'b0000011100111101011100,
    22'b0000011110000101001000,
    22'b0000011111000010100100,
    22'b0000011111100001010010,
    22'b0000011111101011100001,
    22'b0000011111010111000011,
    22'b0000011110100011110110,
    22'b0000011101100110011010,
    22'b0000011100011110101110,
    22'b0000011011100001010010,
    22'b0000011010101110000101,
    22'b0000011010100011110110,
    22'b0000011010101110000101,
    22'b0000011011000010100100,
    22'b0000011011101011100001,
    22'b0000011100101000111101,
    22'b0000011101011100001010,
    22'b0000011110001111010111,
    22'b0000011110111000010100,
    22'b0000011111100001010010,
    22'b0000011111101011100001,
    22'b0000011111101011100001,
    22'b0000011111100001010010,
    22'b0000011111100001010010,
    22'b0000011111110101110001,
    22'b0000100000000000000000,
    22'b0000100000101000111101,
    22'b0000100001000111101100,
    22'b0000100001000111101100,
    22'b0000100001011100001010,
    22'b0000100010001111010111,
    22'b0000100010101110000101,
    22'b0000100010100011110110,
    22'b0000100010100011110110,
    22'b0000100010011001100110,
    22'b0000100010000101001000,
    22'b0000100001110000101001,
    22'b0000100001000111101100,
    22'b0000100000011110101110,
    22'b0000011111110101110001,
    22'b0000011111001100110011,
    22'b0000011110101110000101,
    22'b0000011110100011110110,
    22'b0000011110100011110110,
    22'b0000011110100011110110,
    22'b0000011110100011110110,
    22'b0000011110101110000101,
    22'b0000011111001100110011,
    22'b0000011111101011100001,
    22'b0000011111110101110001,
    22'b0000011111101011100001,
    22'b0000011111101011100001,
    22'b0000011111100001010010,
    22'b0000011111100001010010,
    22'b0000011110101110000101,
    22'b0000011110000101001000,
    22'b0000011101011100001010,
    22'b0000011100010100011111,
    22'b0000011011001100110011,
    22'b0000011010101110000101,
    22'b0000011010101110000101,
    22'b0000011010111000010100,
    22'b0000011011000010100100,
    22'b0000011011100001010010,
    22'b0000011100001010001111,
    22'b0000011100101000111101,
    22'b0000011101000111101100,
    22'b0000100000101000111101,
    22'b0000100001010001111011,
    22'b0000100010001111010111,
    22'b0000100010111000010100,
    22'b0000100010011001100110,
    22'b0000100001111010111000,
    22'b0000100001110000101001,
    22'b0000100001010001111011,
    22'b0000100001011100001010,
    22'b0000100001110000101001,
    22'b0000100001111010111000,
    22'b0000100010001111010111,
    22'b0000100010101110000101,
    22'b0000100011000010100100,
    22'b0000100011010111000011,
    22'b0000100011100001010010,
    22'b0000100011100001010010,
    22'b0000100011001100110011,
    22'b0000100010001111010111,
    22'b0000100001010001111011,
    22'b0000100000010100011111,
    22'b0000011111100001010010,
    22'b0000011111001100110011,
    22'b0000011111000010100100,
    22'b0000011111000010100100,
    22'b0000011111000010100100,
    22'b0000011110100011110110,
    22'b0000011110000101001000,
    22'b0000011101010001111011,
    22'b0000011011101011100001,
    22'b0000011001011100001010,
    22'b0000010110001111010111,
    22'b0000010011101011100001,
    22'b0000010000101000111101,
    22'b0000001101011100001010,
    22'b0000001001110000101001,
    22'b0000000011000010100100,
    22'b1111111111001100110011,
    22'b1111111100011110101110,
    22'b1111111010011001100110,
    22'b1111111001111010111000,
    22'b1111111010101110000101,
    22'b1111111011101011100001,
    22'b1111111011100001010010,
    22'b1111111011001100110011,
    22'b1111111010100011110110,
    22'b1111111001111010111000,
    22'b1111111001011100001010,
    22'b1111111000010100011111,
    22'b1111110111000010100100,
    22'b1111110101111010111000,
    22'b1111110100110011001101,
    22'b1111110100110011001101,
    22'b1111110100111101011100,
    22'b1111110101011100001010,
    22'b1111110110000101001000,
    22'b1111110110100011110110,
    22'b1111110110101110000101,
    22'b1111110111001100110011,
    22'b1111111000000000000000,
    22'b1111111000101000111101,
    22'b1111111001011100001010,
    22'b1111111010000101001000,
    22'b1111111010001111010111,
    22'b1111111010001111010111,
    22'b1111111001111010111000,
    22'b1111111001100110011010,
    22'b1111111001010001111011,
    22'b1111111001010001111011,
    22'b1111111000111101011100,
    22'b1111111000101000111101,
    22'b1111111000010100011111,
    22'b1111110111110101110001,
    22'b1111110111100001010010,
    22'b1111110111000010100100,
    22'b1111110110101110000101,
    22'b1111110110011001100110,
    22'b1111110101111010111000,
    22'b1111110101011100001010,
    22'b1111110100011110101110,
    22'b1111110001011100001010,
    22'b1111101110101110000101,
    22'b1111101100001010001111,
    22'b1111101010001111010111,
    22'b1111101001011100001010,
    22'b1111101110101110000101,
    22'b1111110000011110101110,
    22'b1111110010000101001000,
    22'b1111110011110101110001,
    22'b1111110100111101011100,
    22'b1111110110000101001000,
    22'b1111110111000010100100,
    22'b1111110111110101110001,
    22'b1111111000010100011111,
    22'b1111111000111101011100,
    22'b1111111001011100001010,
    22'b1111111001111010111000,
    22'b1111111010100011110110,
    22'b1111111010101110000101,
    22'b1111111010111000010100,
    22'b1111111010101110000101,
    22'b1111111010100011110110,
    22'b1111111010100011110110,
    22'b1111111010100011110110,
    22'b1111111010011001100110,
    22'b1111111010011001100110,
    22'b1111111010011001100110,
    22'b1111111010001111010111,
    22'b1111111010000101001000,
    22'b1111111001111010111000,
    22'b1111111001100110011010,
    22'b1111111001010001111011,
    22'b1111111000111101011100,
    22'b1111111000011110101110,
    22'b1111111000010100011111,
    22'b1111111000010100011111,
    22'b1111111000010100011111,
    22'b1111111000011110101110,
    22'b1111111000111101011100,
    22'b1111111001000111101100,
    22'b1111111001010001111011,
    22'b1111111001111010111000,
    22'b1111111010000101001000,
    22'b1111111010001111010111,
    22'b1111111000110011001101,
    22'b1111110111110101110001,
    22'b1111110110111000010100,
    22'b1111110101111010111000,
    22'b1111110101010001111011,
    22'b1111110101010001111011,
    22'b1111110101011100001010,
    22'b1111110110000101001000,
    22'b1111110110100011110110,
    22'b1111110110101110000101,
    22'b1111110110101110000101,
    22'b1111110101111010111000,
    22'b1111110100111101011100,
    22'b1111110100000000000000,
    22'b1111110010101110000101,
    22'b1111110001000111101100,
    22'b1111110000001010001111,
    22'b1111101111001100110011,
    22'b1111101110000101001000,
    22'b1111101100110011001101,
    22'b1111101100000000000000,
    22'b1111101011100001010010,
    22'b1111101011010111000011,
    22'b1111101011100001010010,
    22'b1111101011100001010010,
    22'b1111101011010111000011,
    22'b1111101011001100110011,
    22'b1111101010101110000101,
    22'b1111101001111010111000,
    22'b1111100110001111010111,
    22'b1111100101000111101100,
    22'b1111100100011110101110,
    22'b1111100011101011100001,
    22'b1111100011010111000011,
    22'b1111100011000010100100,
    22'b1111100010101110000101,
    22'b1111100010000101001000,
    22'b1111100001011100001010,
    22'b1111100001110000101001,
    22'b1111100010100011110110,
    22'b1111100011010111000011,
    22'b1111100100010100011111,
    22'b1111100101000111101100,
    22'b1111100101100110011010,
    22'b1111100101111010111000,
    22'b1111100110011001100110,
    22'b1111100111000010100100,
    22'b1111101000001010001111,
    22'b1111101001100110011010,
    22'b1111101010100011110110,
    22'b1111101011010111000011,
    22'b1111101011101011100001,
    22'b1111101011001100110011,
    22'b1111101010011001100110,
    22'b1111101001100110011010,
    22'b1111101000000000000000,
    22'b1111101000000000000000,
    22'b1111100111110101110001,
    22'b1111100111101011100001,
    22'b1111100111110101110001,
    22'b1111101000010100011111,
    22'b1111101001011100001010,
    22'b1111101010111000010100,
    22'b1111101011010111000011,
    22'b1111101011110101110001,
    22'b1111101100001010001111,
    22'b1111101100001010001111,
    22'b1111101101000111101100,
    22'b1111101110001111010111,
    22'b1111101110111000010100,
    22'b1111101111110101110001,
    22'b1111110000001010001111,
    22'b1111110000010100011111,
    22'b1111110000110011001101,
    22'b1111110010000101001000,
    22'b1111110010100011110110,
    22'b1111110011100001010010,
    22'b1111110100010100011111,
    22'b1111110100010100011111,
    22'b1111110100011110101110,
    22'b1111110100011110101110,
    22'b1111110100111101011100,
    22'b1111110101011100001010,
    22'b1111110110001111010111,
    22'b1111110111001100110011,
    22'b1111111010000101001000,
    22'b1111111001111010111000,
    22'b1111111001000111101100,
    22'b1111111000010100011111,
    22'b1111110111100001010010,
    22'b1111110110111000010100,
    22'b1111110110100011110110,
    22'b1111110110001111010111,
    22'b1111110101111010111000,
    22'b1111110101010001111011,
    22'b1111110100101000111101,
    22'b1111110100001010001111,
    22'b1111110011101011100001,
    22'b1111110011000010100100,
    22'b1111110010111000010100,
    22'b1111110010101110000101,
    22'b1111110010101110000101,
    22'b1111110010111000010100,
    22'b1111110011000010100100,
    22'b1111110011010111000011,
    22'b1111110011110101110001,
    22'b1111110100010100011111,
    22'b1111110100011110101110,
    22'b1111110100011110101110,
    22'b1111110100010100011111,
    22'b1111110100000000000000,
    22'b1111110011101011100001,
    22'b1111110011001100110011,
    22'b1111110010001111010111,
    22'b1111110001010001111011,
    22'b1111110000011110101110,
    22'b1111101111101011100001,
    22'b1111101110000101001000,
    22'b1111101100111101011100,
    22'b1111101011101011100001,
    22'b1111100100010100011111,
    22'b1111100010111000010100,
    22'b1111100001100110011010,
    22'b1111011111110101110001,
    22'b1111011110111000010100,
    22'b1111011101110000101001,
    22'b1111011101000111101100,
    22'b1111011100101000111101,
    22'b1111011100010100011111,
    22'b1111011100010100011111,
    22'b1111011100011110101110,
    22'b1111011100110011001101,
    22'b1111011101010001111011,
    22'b1111011101111010111000,
    22'b1111011110111000010100,
    22'b1111100000010100011111,
    22'b1111100001011100001010,
    22'b1111100010100011110110,
    22'b1111100011110101110001,
    22'b1111100101011100001010,
    22'b1111100110100011110110,
    22'b1111100111101011100001,
    22'b1111101000111101011100,
    22'b1111101001110000101001,
    22'b1111101010100011110110,
    22'b1111101011001100110011,
    22'b1111101011101011100001,
    22'b1111101011101011100001,
    22'b1111101011101011100001,
    22'b1111101011010111000011,
    22'b1111101010100011110110,
    22'b1111101001100110011010,
    22'b1111101000010100011111,
    22'b1111100110101110000101,
    22'b1111100100001010001111,
    22'b1111100001111010111000,
    22'b1111011111010111000011,
    22'b1111011100010100011111,
    22'b1111011000000000000000,
    22'b1111010100111101011100,
    22'b1111010010101110000101,
    22'b1111010001111010111000,
    22'b1111011000000000000000,
    22'b1111011001111010111000,
    22'b1111011011100001010010,
    22'b1111011101100110011010,
    22'b1111011110111000010100,
    22'b1111100000101000111101,
    22'b1111100010011001100110,
    22'b1111100011110101110001,
    22'b1111100100110011001101,
    22'b1111100101100110011010,
    22'b1111100111000010100100,
    22'b1111101000001010001111,
    22'b1111101000111101011100,
    22'b1111101001110000101001,
    22'b1111101001110000101001,
    22'b1111101001111010111000,
    22'b1111101010100011110110,
    22'b1111101011000010100100,
    22'b1111101010111000010100,
    22'b1111101011000010100100,
    22'b1111101010111000010100,
    22'b1111101001100110011010,
    22'b1111100110111000010100,
    22'b1111100100010100011111,
    22'b1111100001010001111011,
    22'b1111011100010100011111,
    22'b1111010100001010001111,
    22'b1111001110000101001000,
    22'b1111000111001100110011,
    22'b1111000001111010111000,
    22'b1110111110101110000101,
    22'b1110111011110101110001,
    22'b1110111000111101011100,
    22'b1110110110000101001000,
    22'b1110110011110101110001,
    22'b1110110010101110000101,
    22'b1110110010000101001000,
    22'b1110110110101110000101,
    22'b1110111101110000101001,
    22'b1111010000101000111101,
    22'b1111010011000010100100,
    22'b1111010100011110101110,
    22'b1111010110101110000101,
    22'b1111010111100001010010,
    22'b1111011000101000111101,
    22'b1111011001111010111000,
    22'b1111011011000010100100,
    22'b1111011101010001111011,
    22'b1111011110100011110110,
    22'b1111011111000010100100,
    22'b1111011111110101110001,
    22'b1111100000101000111101,
    22'b1111100001011100001010,
    22'b1111100010011001100110,
    22'b1111100011101011100001,
    22'b1111100100000000000000,
    22'b1111100100000000000000,
    22'b1111100100001010001111,
    22'b1111100011001100110011,
    22'b1111100001111010111000,
    22'b1111100000001010001111,
    22'b1111011110101110000101,
    22'b1111011100010100011111,
    22'b1111011010101110000101,
    22'b1111011000010100011111,
    22'b1111010110011001100110,
    22'b1111010011100001010010,
    22'b1111010001000111101100,
    22'b1111010000010100011111,
    22'b1111001100101000111101,
    22'b1111001010000101001000,
    22'b1111001010111000010100,
    22'b1111001000111101011100,
    22'b1111010101011100001010,
    22'b1111011101000111101100,
    22'b1111100010101110000101,
    22'b1111101000011110101110,
    22'b1111101011010111000011,
    22'b1111101101011100001010,
    22'b1111101111010111000011,
    22'b1111110000110011001101,
    22'b1111110001100110011010,
    22'b1111110001110000101001,
    22'b1111110001000111101100,
    22'b1111110000011110101110,
    22'b1111110000011110101110,
    22'b1111110001000111101100,
    22'b1111110010000101001000,
    22'b1111110011010111000011,
    22'b1111110100001010001111,
    22'b1111110100101000111101,
    22'b1111110101000111101100,
    22'b1111110100111101011100,
    22'b1111110100111101011100,
    22'b1111110101010001111011,
    22'b1111110101000111101100,
    22'b1111110100111101011100,
    22'b1111110100010100011111,
    22'b1111110100001010001111,
    22'b1111110011100001010010,
    22'b1111110010000101001000,
    22'b1111110001111010111000,
    22'b1111110001110000101001,
    22'b1111110011000010100100,
    22'b1111110100000000000000,
    22'b1111110100001010001111,
    22'b1111110100001010001111,
    22'b1111110000011110101110,
    22'b1111110000000000000000,
    22'b1111101111010111000011,
    22'b1111101111000010100100,
    22'b1111101110101110000101,
    22'b1111101111010111000011,
    22'b1111110000000000000000,
    22'b1111110000011110101110,
    22'b1111101111100001010010,
    22'b1111101110000101001000,
    22'b1111101101010001111011,
    22'b1111101100101000111101,
    22'b1111101011010111000011,
    22'b1111101001110000101001,
    22'b1111101000011110101110,
    22'b1111100111000010100100,
    22'b1111100101000111101100,
    22'b1111100010101110000101,
    22'b1111011110011001100110,
    22'b1111010111110101110001,
    22'b1111010010100011110110,
    22'b1111001100000000000000,
    22'b1111001000011110101110,
    22'b1111000100110011001101,
    22'b1111000001011100001010,
    22'b1110111111000010100100,
    22'b1110111100101000111101,
    22'b1110111010111000010100,
    22'b1110111001100110011010,
    22'b1110111000010100011111,
    22'b1110111000000000000000,
    22'b1110111000101000111101,
    22'b1110111010000101001000,
    22'b1110111100110011001101,
    22'b1111000000011110101110,
    22'b1111000110111000010100,
    22'b1111010101000111101100,
    22'b1111010101111010111000,
    22'b1111010110101110000101,
    22'b1111010111001100110011,
    22'b1111010111010111000011,
    22'b1111010111001100110011,
    22'b1111010101111010111000,
    22'b1111010100111101011100,
    22'b1111010011101011100001,
    22'b1111010001110000101001,
    22'b1111010000101000111101,
    22'b1111001111110101110001,
    22'b1111001111101011100001,
    22'b1111001111001100110011,
    22'b1111001111001100110011,
    22'b1111001111000010100100,
    22'b1111001111010111000011,
    22'b1111010000001010001111,
    22'b1111010000111101011100,
    22'b1111010001110000101001,
    22'b1111010011000010100100,
    22'b1111010100001010001111,
    22'b1111010101110000101001,
    22'b1111010111110101110001,
    22'b1111011011100001010010,
    22'b1111011110011001100110,
    22'b1111100000111101011100,
    22'b1111100011010111000011,
    22'b1111100101111010111000,
    22'b1111100111100001010010,
    22'b1111101000111101011100,
    22'b1111101010011001100110,
    22'b1111101010101110000101,
    22'b1111101010001111010111,
    22'b1111101001111010111000,
    22'b1111101010001111010111,
    22'b1111101010111000010100,
    22'b1111101011100001010010,
    22'b1111101100111101011100,
    22'b1111101110011001100110,
    22'b1111110000001010001111,
    22'b1111110001111010111000,
    22'b1111110100010100011111,
    22'b1111110101011100001010,
    22'b1111110110000101001000,
    22'b1111110101110000101001,
    22'b1111110100111101011100,
    22'b1111110011110101110001,
    22'b1111110010101110000101,
    22'b1111110001000111101100,
    22'b1111101111110101110001,
    22'b1111101110101110000101,
    22'b1111101101111010111000,
    22'b1111101101111010111000,
    22'b1111101110100011110110,
    22'b1111101111110101110001,
    22'b1111110000110011001101,
    22'b1111110010011001100110,
    22'b1111110100110011001101,
    22'b1111111000000000000000,
    22'b1111111010101110000101,
    22'b1111111101110000101001,
    22'b0000000001110000101001,
    22'b0000001101010001111011,
    22'b0000001101100110011010,
    22'b0000001100111101011100,
    22'b0000001011100001010010,
    22'b0000001000010100011111,
    22'b0000000101011100001010,
    22'b0000000010001111010111,
    22'b1111111101011100001010,
    22'b1111111000111101011100,
    22'b1111110101000111101100,
    22'b1111110010100011110110,
    22'b1111101111100001010010,
    22'b1111101101111010111000,
    22'b1111101100111101011100,
    22'b1111101100001010001111,
    22'b1111101100001010001111,
    22'b1111101100110011001101,
    22'b1111101101010001111011,
    22'b1111101101011100001010,
    22'b1111101101011100001010,
    22'b1111101101000111101100,
    22'b1111101011100001010010,
    22'b1111101000011110101110,
    22'b1111100111010111000011,
    22'b1111100111101011100001,
    22'b1111100111100001010010,
    22'b1111101001100110011010,
    22'b1111101100101000111101,
    22'b1111101111100001010010,
    22'b1111110011100001010010,
    22'b1111110110111000010100,
    22'b1111111011101011100001,
    22'b1111111011000010100100,
    22'b1111111010100011110110,
    22'b1111111001111010111000,
    22'b1111111001011100001010,
    22'b1111111001010001111011,
    22'b1111111001000111101100,
    22'b1111111000111101011100,
    22'b1111111000111101011100,
    22'b1111111001000111101100,
    22'b1111111000111101011100,
    22'b1111111000101000111101,
    22'b1111110111101011100001,
    22'b1111110110100011110110,
    22'b1111110101100110011010,
    22'b1111110100110011001101,
    22'b1111110011110101110001,
    22'b1111110011010111000011,
    22'b1111110010111000010100,
    22'b1111110010011001100110,
    22'b1111110010001111010111,
    22'b1111110010001111010111,
    22'b1111110010100011110110,
    22'b1111110011000010100100,
    22'b1111110111100001010010,
    22'b1111111000101000111101,
    22'b1111111001111010111000,
    22'b1111111010101110000101,
    22'b1111111011001100110011,
    22'b1111111011101011100001,
    22'b1111111100001010001111,
    22'b1111111100011110101110,
    22'b1111111100110011001101,
    22'b1111111101000111101100,
    22'b1111111101010001111011,
    22'b1111111101011100001010,
    22'b1111111101011100001010,
    22'b1111111101010001111011,
    22'b1111111101010001111011,
    22'b1111111101000111101100,
    22'b1111111100111101011100,
    22'b1111111100011110101110,
    22'b1111111100010100011111,
    22'b1111111100010100011111,
    22'b1111111100010100011111,
    22'b1111111100101000111101,
    22'b1111111101000111101100,
    22'b1111111101100110011010,
    22'b1111111110011001100110,
    22'b0000000000101000111101,
    22'b0000000000111101011100,
    22'b0000000001100110011010,
    22'b0000000010000101001000,
    22'b0000000010111000010100,
    22'b0000000011101011100001,
    22'b0000000100110011001101,
    22'b0000000101011100001010,
    22'b0000000110001111010111,
    22'b0000000111000010100100,
    22'b0000001000001010001111,
    22'b0000001001000111101100,
    22'b0000001010000101001000,
    22'b0000001011001100110011,
    22'b0000001100110011001101,
    22'b0000001110000101001000,
    22'b0000001111000010100100,
    22'b0000001111110101110001,
    22'b0000001100101000111101,
    22'b0000001001111010111000,
    22'b0000000111101011100001,
    22'b0000000011110101110001,
    22'b1111111111001100110011,
    22'b1111111011110101110001,
    22'b1111111001100110011010,
    22'b1111111001010001111011,
    22'b1111111001110000101001,
    22'b1111111011001100110011,
    22'b1111111100110011001101,
    22'b1111111110000101001000,
    22'b1111111111000010100100,
    22'b1111111111100001010010,
    22'b0000000010001111010111,
    22'b0000000001110000101001,
    22'b0000000001011100001010,
    22'b0000000000111101011100,
    22'b1111111111110101110001,
    22'b1111111101100110011010,
    22'b1111111100101000111101,
    22'b1111111100000000000000,
    22'b1111111010100011110110,
    22'b1111111000110011001101,
    22'b1111111000001010001111,
    22'b1111110111110101110001,
    22'b1111111000000000000000,
    22'b1111111000001010001111,
    22'b1111111000101000111101,
    22'b1111111001010001111011,
    22'b1111111010000101001000,
    22'b1111111010111000010100,
    22'b1111111011010111000011,
    22'b1111111011010111000011,
    22'b1111111011001100110011,
    22'b1111111010111000010100,
    22'b1111111010001111010111,
    22'b1111111001111010111000,
    22'b1111111001100110011010,
    22'b1111111010001111010111,
    22'b1111111010111000010100,
    22'b1111111011001100110011,
    22'b1111111010101110000101,
    22'b1111111010001111010111,
    22'b1111111001011100001010,
    22'b1111110100111101011100,
    22'b1111110101100110011010,
    22'b1111110101011100001010,
    22'b1111110100110011001101,
    22'b1111110100010100011111,
    22'b1111110100000000000000,
    22'b1111110011100001010010,
    22'b1111110011000010100100,
    22'b1111110010001111010111,
    22'b1111110001111010111000,
    22'b1111110001111010111000,
    22'b1111110010000101001000,
    22'b1111110010011001100110,
    22'b1111110010101110000101,
    22'b1111110011001100110011,
    22'b1111110100000000000000,
    22'b1111110100011110101110,
    22'b1111110100110011001101,
    22'b1111110100110011001101,
    22'b1111110100101000111101,
    22'b1111110100010100011111,
    22'b1111110011101011100001,
    22'b1111110010111000010100,
    22'b1111110001000111101100,
    22'b1111110000111101011100,
    22'b1111110000110011001101,
    22'b1111110000110011001101,
    22'b1111110000110011001101,
    22'b1111110000101000111101,
    22'b1111110000110011001101,
    22'b1111110000110011001101,
    22'b1111110000111101011100,
    22'b1111110001100110011010,
    22'b1111110001000111101100,
    22'b1111110000110011001101,
    22'b1111110000001010001111,
    22'b1111101111001100110011,
    22'b1111101101111010111000,
    22'b1111101101010001111011,
    22'b1111101100001010001111,
    22'b1111101010101110000101,
    22'b1111101001011100001010,
    22'b1111100111010111000011,
    22'b1111100100101000111101,
    22'b1111100000101000111101,
    22'b1111011101010001111011,
    22'b1111011001111010111000,
    22'b1111010110111000010100,
    22'b1111010100000000000000,
    22'b1111010010111000010100,
    22'b1111010101010001111011,
    22'b1111010101110000101001,
    22'b1111010110101110000101,
    22'b1111010101111010111000,
    22'b1111010101000111101100,
    22'b1111010101011100001010,
    22'b1111010110111000010100,
    22'b1111011001010001111011,
    22'b1111100011010111000011,
    22'b1111101001011100001010,
    22'b1111101101010001111011,
    22'b1111110011001100110011,
    22'b1111111010111000010100,
    22'b1111111110101110000101,
    22'b0000000000111101011100,
    22'b0000000010011001100110,
    22'b0000000011101011100001,
    22'b0000000011110101110001,
    22'b0000000010101110000101,
    22'b0000000001110000101001,
    22'b0000000010101110000101,
    22'b0000000010011001100110,
    22'b0000000001110000101001,
    22'b0000000001111010111000,
    22'b0000000001011100001010,
    22'b0000000000101000111101,
    22'b0000000000010100011111,
    22'b0000000000000000000000,
    22'b1111111110111000010100,
    22'b1111111101100110011010,
    22'b1111111100101000111101,
    22'b1111111011101011100001,
    22'b1111111010000101001000,
    22'b1111111000110011001101,
    22'b1111110100000000000000,
    22'b1111110011100001010010,
    22'b1111110011010111000011,
    22'b1111110011100001010010,
    22'b1111110100000000000000,
    22'b1111110101010001111011,
    22'b1111110110100011110110,
    22'b1111110111101011100001,
    22'b1111111010000101001000,
    22'b1111111100011110101110,
    22'b1111111111000010100100,
    22'b0000000001110000101001,
    22'b0000000101110000101001,
    22'b0000001000010100011111,
    22'b0000001010101110000101,
    22'b0000001100110011001101,
    22'b0000001111000010100100,
    22'b0000010000001010001111,
    22'b0000010000101000111101,
    22'b0000010000011110101110,
    22'b0000010000000000000000,
    22'b0000001111101011100001,
    22'b0000001111001100110011,
    22'b0000001111000010100100,
    22'b0000001111001100110011,
    22'b0000001111101011100001,
    22'b0000010000010100011111,
    22'b0000010001110000101001,
    22'b0000010010111000010100,
    22'b0000010011100001010010,
    22'b0000010100000000000000,
    22'b0000010100101000111101,
    22'b0000010101000111101100,
    22'b0000010101011100001010,
    22'b0000010101100110011010,
    22'b0000010101010001111011,
    22'b0000010100011110101110,
    22'b0000010011010111000011,
    22'b0000001011110101110001,
    22'b0000001010101110000101,
    22'b0000001010011001100110,
    22'b0000001010111000010100,
    22'b0000001100110011001101,
    22'b0000001111000010100100,
    22'b0000010001000111101100,
    22'b0000010011110101110001,
    22'b0000010111001100110011,
    22'b0000011000110011001101,
    22'b0000011001111010111000,
    22'b0000011010011001100110,
    22'b0000011010001111010111,
    22'b0000011001110000101001,
    22'b0000011000110011001101,
    22'b0000010111101011100001,
    22'b0000010101100110011010,
    22'b0000010100001010001111,
    22'b0000010011100001010010,
    22'b0000010011001100110011,
    22'b0000010011110101110001,
    22'b0000010100101000111101,
    22'b0000010101110000101001,
    22'b0000010111100001010010,
    22'b0000011000110011001101,
    22'b0000011001011100001010,
    22'b0000011001110000101001,
    22'b0000011011100001010010,
    22'b0000011100111101011100,
    22'b0000011110111000010100,
    22'b0000100000011110101110,
    22'b0000100010000101001000,
    22'b0000100010100011110110,
    22'b0000100010011001100110,
    22'b0000100001111010111000,
    22'b0000100000110011001101,
    22'b0000011111110101110001,
    22'b0000011111001100110011,
    22'b0000011110101110000101,
    22'b0000011110101110000101,
    22'b0000011111000010100100,
    22'b0000011111110101110001,
    22'b0000100110001111010111,
    22'b0000100111100001010010,
    22'b0000101000101000111101,
    22'b0000101001011100001010,
    22'b0000101010111000010100,
    22'b0000101100000000000000,
    22'b0000101101011100001010,
    22'b0000101110111000010100,
    22'b0000110000111101011100,
    22'b0000110010111000010100,
    22'b0000110101000111101100,
    22'b0000110111110101110001,
    22'b0000111011010111000011,
    22'b0000111101011100001010,
    22'b0000111111001100110011,
    22'b0001000000011110101110,
    22'b0001000001011100001010,
    22'b0001000001010001111011,
    22'b0001000000010100011111,
    22'b0000111110111000010100,
    22'b0000111100111101011100,
    22'b0000111011010111000011,
    22'b0000111001111010111000,
    22'b0000111000011110101110,
    22'b0000110110111000010100,
    22'b0000110110000101001000,
    22'b0000110101100110011010,
    22'b0000110101011100001010,
    22'b0000110101011100001010,
    22'b0000110101011100001010,
    22'b0000110101011100001010,
    22'b0000110101010001111011,
    22'b0000110100110011001101,
    22'b0000110100010100011111,
    22'b0000110011101011100001,
    22'b0000110010111000010100,
    22'b0000110010001111010111,
    22'b0000110001010001111011,
    22'b0000110000101000111101,
    22'b0000101111110101110001,
    22'b0000101111001100110011,
    22'b0000101110001111010111,
    22'b0000101101011100001010,
    22'b0000101100111101011100,
    22'b0000101100010100011111,
    22'b0000101011110101110001,
    22'b0000101011001100110011,
    22'b0000101010011001100110,
    22'b0000101001011100001010,
    22'b0000101000010100011111,
    22'b0000100110100011110110,
    22'b0000100101000111101100,
    22'b0000100011101011100001,
    22'b0000100010011001100110,
    22'b0000100000110011001101,
    22'b0000011111100001010010,
    22'b0000011110001111010111,
    22'b0000011101000111101100,
    22'b0000011100001010001111,
    22'b0000011011101011100001,
    22'b0000011100000000000000,
    22'b0000011100011110101110,
    22'b0000011101000111101100,
    22'b0000011101110000101001,
    22'b0000011110000101001000,
    22'b0000011110011001100110
};

